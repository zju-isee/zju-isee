// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Fri Jun 09 10:06:12 2023
//
// Verilog Description of module LED
//

module LED (clk_50m, reset_n, led_col, led_row) /* synthesis syn_module_defined=1 */ ;   // led.v(1[8:11])
    input clk_50m;   // led.v(3[11:18])
    input reset_n;   // led.v(3[19:26])
    output [7:0]led_col;   // led.v(4[18:25])
    output [7:0]led_row;   // led.v(5[18:25])
    
    wire clk_50m_c /* synthesis SET_AS_NETWORK=clk_50m_c, is_clock=1 */ ;   // led.v(3[11:18])
    
    wire reset_n_c;
    wire [15:0]cnt_scan;   // led.v(7[16:24])
    
    wire led_row_c_7, led_row_c_6, led_row_c_5, led_row_c_4, led_row_c_3, 
        led_row_c_2, led_row_c_1, led_row_c_0;
    wire [7:0]col_buf;   // led.v(8[23:30])
    wire [25:0]cnt_next;   // led.v(9[16:24])
    wire [6:0]scan_data;   // led.v(10[15:24])
    
    wire n78, n76, n1679, n2770;
    wire [7:0]col3;   // led.v(11[25:29])
    
    wire n81;
    wire [7:0]col4;   // led.v(11[30:34])
    
    wire n3228, n844, n3167, n789, n73, n2466, n2586, n1582, 
        n3225, n3165, n3163, n3161, n824, n3196, n3193, n3190, 
        n3187, n3184, n3181, n3178, n3175, n70, n817, n3231, 
        n70_adj_1, n776, n81_adj_2, n2752, n836, n2423, n64, n48, 
        n3200, n73_adj_3, n3203, n2758, n78_adj_4, n829, n2760, 
        n775, n819, n3234, n2784, n3206, n67, n28, n3159, n841, 
        n661, n814, n790, n81_adj_5, n787, n14, n3212, n3215, 
        n76_adj_6, n78_adj_7, n2764, n39, n6, n37, n32, n3222, 
        n67_adj_8, n3219, n70_adj_9, n786, n81_adj_10, n10, n27, 
        n3209, n76_adj_11, n78_adj_12, n3197, n26, col1_7__N_71, 
        col1_7__N_72, col1_7__N_74, n2593, n3363, n8, n813, n831, 
        n2757, n785, n465, n788, n81_adj_13, n3152, n818, n835, 
        n2789, n845, n1580, n3157, n78_adj_14, n73_adj_15, n3237, 
        n812, n8_adj_16, n773, n81_adj_17, n3150, n792, n816, 
        n1588, n67_adj_18, n3246, n78_adj_19, n76_adj_20, n3240, 
        n73_adj_21, n3243, n784, n828, n3153, n81_adj_22, n791, 
        n815, n67_adj_23, n3255, n78_adj_24, n76_adj_25, n3252, 
        n10_adj_26, n3249, n820, n832, n33, n3258, n27_adj_27, 
        n6_adj_28, n19, n30, n32_adj_29, n847, n3261, n29, n27_adj_30, 
        n24, n30_adj_31, n32_adj_32, n30_adj_33, n4, n3264, n11, 
        n15, n18, n29_adj_34, n27_adj_35, n22, n1574, n2494, n2407, 
        n30_adj_36, n3267, n28_adj_37, n27_adj_38, n2628, n28_adj_39, 
        n3270, n30_adj_40, n14_adj_41, n7, n14_adj_42, n1578, n14_adj_43, 
        n3276, n846, n1572, n3173, n20, n23, n21, n3285, n18_adj_44, 
        n14_adj_45, n157, n84, n156, n155, n154, n153, n151, 
        n150, n149, n148, n147, n75, n146, n145, n144, n143, 
        n142, n141, n140, n139, n138, n137, n136, n2579, n23_adj_46, 
        n3288, n135, n134, n130, n129, n128, n133, n28_adj_47, 
        n27_adj_48, n3291, n126, n125, n124, n123, n122, n121, 
        n3294, n120, n119, n118, n117, n21_adj_49, n3297, n116, 
        n115, n114, n113, n112, n111, n110, n109, n108, n2773, 
        n3300, n106, n83, n107, n2614, n25, n726, n3303, n6_adj_50, 
        n1656, n2557, n3306, n2777, n1628, n79, n3309, n2550, 
        n3312, n3315, n1624, n127, n152, n2437, pwr, n15_adj_51, 
        n22_adj_52, n18_adj_53, n3318, n4_adj_54, n5, n3321, n78_adj_55, 
        n85, n2733, n2726, n3324, n12, n34, n31, n2719, n1727, 
        n1622, n2712, n2754, n659, n3330, n5_adj_56, n3327, n21_adj_57, 
        n23_adj_58, n2705, n3333, n2698, n20_adj_59, n2691, n3210, 
        n39_adj_60, n38, n2430, n25_adj_61, n37_adj_62, n36, n35, 
        n34_adj_63, n2508, n3345, n3351, n3348, n82, n3357, n1618, 
        n3360, n81_adj_64, n7_adj_65, n49, n7_adj_66, n4_adj_67, 
        n70_adj_68, n5_adj_69, n10_adj_70, n12_adj_71, n8_adj_72, 
        n2543, n8_adj_73, n1719, n6_adj_74, n20_adj_75, n3273, n4_adj_76, 
        n3279, n3365, n3364, n805, n3342, n19_adj_77, n3339, n2684, 
        n2536, n18_adj_78, n2416, n3336, n2677, n71, n72, n3362, 
        n73_adj_79, n74, n3354, n76_adj_80, n780, n77, n2748, 
        n80, n3361, n3359, n3358, n3356, n1614, n1717, n3355, 
        n2515, n4_adj_81, n3353, n3156, n1709, n2670, n2501, n2663, 
        n3151, n3352, n3350, n3349, n2529, n3347, n2656, n1576, 
        n1586, n3346, n1606, n3343, n3341, n1699, n1695, n3340, 
        n3338, n2778, n3337, n3335, n1685, n3334, n3332, n1681, 
        n2649, n3331, gnd, n2522, n2642, n28_adj_82, n3329, n3328, 
        n3326, n27_adj_83, n26_adj_84, n3325, n2444, n3323, n2635, 
        n24_adj_85, n3322, n2473, n5_adj_86, n3320, n2621, n2480, 
        n2607, n3319, n3317, n3316, n2487, n23_adj_87, n3314, 
        n2600, n3313, n3311, n3310, n3308, n22_adj_88, n21_adj_89, 
        n3307, n14_adj_90, n13, n20_adj_91, n3305, n3304, n3302, 
        n3301, n3299, n3298, n3296, n3295, n3293, n3292, n3290, 
        n3289, n3287, n3286, n3284, n3283, n3282, n3280, n3278, 
        n3277, n19_adj_92, n3275, n3274, n3272, n3271, n3269, 
        n3268, n3265, n18_adj_93, n3263, n3262, n3260, n3259, 
        n3257, n3256, n3254, n3253, n3251, n3250, n3248, n3247, 
        n3245, n3244, n3242, n3241, n3239, n3238, n3236, n3235, 
        n3233, n3232, n3230, n3229, n3227, n3226, n3224, n3223, 
        n4_adj_94, n3221, n3220, n3218, n3217, n3216, n3214, n3213, 
        n3211, n3208, n3194, n3207, n3191, n3205, n3188, n3204, 
        n3185, n3202, n3182, n3201, n3179, n12_adj_95, n19_adj_96, 
        n3199, n3176, n3198, n12_adj_97, n28_adj_98, n3171;
    
    AND2 i2311 (.O(n2642), .I0(n2635), .I1(cnt_next[10]));
    DFFCS row_buf_i0_i8 (.Q(led_row_c_7), .D(led_row_c_6), .CLK(clk_50m_c), 
          .CE(n847), .S(reset_n_c));   // led.v(26[13] 35[11])
    OR2 i2875 (.O(n3202), .I0(n3201), .I1(n3200));
    AND2 i2318 (.O(n2649), .I0(n2642), .I1(cnt_next[11]));
    OR2 i1 (.O(n81_adj_13), .I0(n2752), .I1(n73_adj_15));
    OR2 i1_adj_1 (.O(n78_adj_14), .I0(n2754), .I1(n3151));
    AND2 i2325 (.O(n2656), .I0(n2649), .I1(cnt_next[12]));
    AND2 i2099 (.O(n2430), .I0(n2423), .I1(scan_data[3]));
    OR3 i2 (.O(n2777), .I0(n14_adj_43), .I1(scan_data[2]), .I2(scan_data[3]));
    OR2 i2842 (.O(n3171), .I0(n1580), .I1(n1695));
    OR2 i2830 (.O(n3159), .I0(n1582), .I1(n1606));
    OR3 i2847 (.O(col_buf[0]), .I0(n1580), .I1(n3173), .I2(led_row_c_4));
    AND2 i2850 (.O(col_buf[1]), .I0(n3176), .I1(n3175));
    AND2 i1_adj_2 (.O(n790), .I0(n784), .I1(n78_adj_19));
    XOR2 i31 (.O(n19_adj_96), .I0(scan_data[2]), .I1(n6_adj_50));
    AND2 i1_adj_3 (.O(n3151), .I0(n3150), .I1(n3272));
    AND4 i2907 (.O(n3234), .I0(led_row_c_4), .I1(n792), .I2(n2784), 
         .I3(n3302));
    OR2 i1_adj_4 (.O(n12_adj_95), .I0(n19_adj_96), .I1(n25));
    AND2 i2853 (.O(col_buf[2]), .I0(n3179), .I1(n3178));
    AND2 i2856 (.O(col_buf[3]), .I0(n3182), .I1(n3181));
    AND2 i1_adj_5 (.O(n791), .I0(n784), .I1(n78_adj_14));
    AND2 i2859 (.O(col_buf[4]), .I0(n3185), .I1(n3184));
    OR3 i2_adj_6 (.O(n2773), .I0(scan_data[0]), .I1(n8_adj_73), .I2(n12_adj_71));
    AND2 i2862 (.O(col_buf[5]), .I0(n3188), .I1(n3187));
    AND2 i7 (.O(n23_adj_46), .I0(cnt_scan[14]), .I1(cnt_scan[11]));
    AND3 i2877 (.O(n3204), .I0(n841), .I1(led_row_c_1), .I2(n30_adj_36));
    AND2 i2865 (.O(col_buf[6]), .I0(n3191), .I1(n3190));
    AND2 i2868 (.O(col_buf[7]), .I0(n3194), .I1(n3193));
    AND2 i2332 (.O(n2663), .I0(n2656), .I1(cnt_next[13]));
    AND6 i15 (.O(n847), .I0(n28_adj_98), .I1(cnt_scan[6]), .I2(n18_adj_78), 
         .I3(n26), .I4(n27), .I5(cnt_scan[0]));
    VCC i2845 (.X(pwr));
    OR2 i1_adj_7 (.O(n81), .I0(n2757), .I1(n2758));
    OR2 i1_adj_8 (.O(n78_adj_4), .I0(n70), .I1(n3153));
    AND4 i2904 (.O(n3231), .I0(led_row_c_2), .I1(n824), .I2(n3215), 
         .I3(n14_adj_45));
    AND3 i2901 (.O(n3228), .I0(col3[3]), .I1(n3215), .I2(led_row_c_2));
    AND3 i2898 (.O(n3225), .I0(col3[3]), .I1(n2784), .I2(led_row_c_4));
    OR2 i1251 (.O(n1588), .I0(led_row_c_0), .I1(led_row_c_1));
    OR2 i2878 (.O(n3205), .I0(n3204), .I1(n3203));
    AND3 i2_adj_9 (.O(n6), .I0(n2789), .I1(n3214), .I2(n39));
    OR2 i1_adj_10 (.O(n81_adj_2), .I0(n76), .I1(n73));
    AND4 i2896 (.O(n3223), .I0(n10), .I1(n824), .I2(led_row_c_7), .I3(n27_adj_27));
    OR2 i2897 (.O(n3224), .I0(n3223), .I1(n3222));
    AND3 i2899 (.O(n3226), .I0(n4_adj_94), .I1(led_row_c_5), .I2(n3311));
    AND3 i2_adj_11 (.O(n2754), .I0(n7_adj_65), .I1(n3278), .I2(n820));
    OR2 i1_adj_12 (.O(n78), .I0(n70_adj_1), .I1(n3152));
    OR2 i1241 (.O(n1578), .I0(n846), .I1(led_row_c_2));
    OR2 i2900 (.O(n3227), .I0(n3226), .I1(n3225));
    AND4 i2895 (.O(n3222), .I0(led_row_c_6), .I1(n805), .I2(n2789), 
         .I3(n3332));
    AND2 i2902 (.O(n3229), .I0(led_row_c_3), .I1(n775));
    INV i1240 (.O(n48), .I0(n1576));
    OR2 i2903 (.O(n3230), .I0(n3229), .I1(n3228));
    AND2 i2892 (.O(n3219), .I0(n14), .I1(n8_adj_16));
    AND3 i2905 (.O(n3232), .I0(n3287), .I1(led_row_c_3), .I2(n773));
    OR2 i2906 (.O(n3233), .I0(n3232), .I1(n3231));
    INV i1363 (.O(n841), .I0(n1699));
    AND4 i2908 (.O(n3235), .I0(n6_adj_28), .I1(n15_adj_51), .I2(led_row_c_5), 
         .I3(n5_adj_56));
    AND2 i2339 (.O(n2670), .I0(n2663), .I1(cnt_next[14]));
    OR2 i2909 (.O(n3236), .I0(n3235), .I1(n3234));
    AND2 i2911 (.O(n3238), .I0(led_row_c_7), .I1(n64));
    AND2 i8 (.O(n24), .I0(cnt_scan[15]), .I1(cnt_scan[9]));
    INV i1361 (.O(n726), .I0(n2777));
    AND2 i2880 (.O(n3207), .I0(led_row_c_7), .I1(n64));
    OR2 i2912 (.O(n3239), .I0(n3238), .I1(n3237));
    AND4 i2914 (.O(n3241), .I0(n22), .I1(n1628), .I2(led_row_c_5), .I3(n5_adj_86));
    AND2 i2_adj_13 (.O(n67_adj_23), .I0(n8), .I1(n3254));
    AND2 i2_adj_14 (.O(n76_adj_25), .I0(n7_adj_66), .I1(n3251));
    OR2 i2915 (.O(n3242), .I0(n3241), .I1(n3240));
    OR2 i1243 (.O(n1580), .I0(led_row_c_2), .I1(led_row_c_3));
    AND3 i2917 (.O(n3244), .I0(n841), .I1(led_row_c_1), .I2(n14_adj_42));
    AND2 i2_adj_15 (.O(n30_adj_31), .I0(n7), .I1(n29));
    OR2 i2832 (.O(n3161), .I0(led_row_c_4), .I1(n3156));
    INV i1359 (.O(n792), .I0(n1695));
    OR2 i2918 (.O(n3245), .I0(n3244), .I1(n3243));
    OR2 i1235 (.O(n1572), .I0(scan_data[3]), .I1(scan_data[4]));
    AND3 i2920 (.O(n3247), .I0(n3308), .I1(led_row_c_5), .I2(n28));
    OR2 i2921 (.O(n3248), .I0(n3247), .I1(n3246));
    INV i1383 (.O(n10_adj_70), .I0(n1719));
    AND2 i2923 (.O(n3250), .I0(led_row_c_7), .I1(n64));
    AND2 i2_adj_16 (.O(n18_adj_44), .I0(n4_adj_67), .I1(scan_data[0]));
    OR2 i2924 (.O(n3251), .I0(n3250), .I1(n3249));
    AND4 i2926 (.O(n3253), .I0(n39), .I1(n824), .I2(led_row_c_1), .I3(n14_adj_43));
    OR2 i2927 (.O(n3254), .I0(n3253), .I1(n3252));
    INV i1381 (.O(n773), .I0(n1717));
    AND2 i2076 (.O(n2407), .I0(scan_data[0]), .I1(n465));
    OR2 i1237 (.O(n1574), .I0(n845), .I1(led_row_c_6));
    OR2 i1_adj_17 (.O(n844), .I0(n12_adj_71), .I1(n11));
    AND2 i2929 (.O(n3256), .I0(scan_data[2]), .I1(n19));
    AND2 i1_adj_18 (.O(n19), .I0(n11), .I1(scan_data[1]));
    OR2 i2930 (.O(n3257), .I0(n3256), .I1(n3255));
    AND2 i2346 (.O(n2677), .I0(n2670), .I1(cnt_next[15]));
    AND2 i2932 (.O(n3259), .I0(scan_data[2]), .I1(scan_data[1]));
    OR2 i2834 (.O(n3163), .I0(led_row_c_0), .I1(n1695));
    OR2 i2933 (.O(n3260), .I0(n3259), .I1(n3258));
    AND2 i2935 (.O(n3262), .I0(scan_data[2]), .I1(n19));
    OR2 i2936 (.O(n3263), .I0(n3262), .I1(n3261));
    AND2 i2885 (.O(n3212), .I0(n10), .I1(n3211));
    AND2 i2297 (.O(n2628), .I0(n2621), .I1(cnt_next[8]));
    AND2 i2353 (.O(n2684), .I0(n2677), .I1(cnt_next[16]));
    AND2 i10 (.O(n26), .I0(n20_adj_75), .I1(n19_adj_77));
    AND2 i11 (.O(n27), .I0(n22_adj_52), .I1(n21_adj_57));
    INV i1238 (.O(n64), .I0(n1574));
    INV i2831 (.O(n4_adj_81), .I0(n3159));
    OR2 i2836 (.O(n3165), .I0(n1695), .I1(n20));
    OR2 i1_adj_19 (.O(n78_adj_12), .I0(n2770), .I1(n67));
    INV i2460 (.O(n2789), .I0(led_row_c_7));
    AND2 i2360 (.O(n2691), .I0(n2684), .I1(cnt_next[17]));
    DFFR cnt_scan_155__i0 (.Q(cnt_scan[0]), .D(n85), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(28[23:33])
    OR2 i1_adj_20 (.O(n81_adj_5), .I0(n76_adj_11), .I1(n2764));
    OR2 i2881 (.O(n3208), .I0(n3207), .I1(n3206));
    AND2 i2938 (.O(n3265), .I0(scan_data[1]), .I1(n11));
    OR2 i1245 (.O(n1582), .I0(led_row_c_4), .I1(led_row_c_5));
    AND3 i2882 (.O(n3209), .I0(col1_7__N_72), .I1(n2784), .I2(led_row_c_1));
    XOR2 i325 (.O(n661), .I0(led_row_c_5), .I1(led_row_c_4));
    AND2 i2941 (.O(n3268), .I0(scan_data[0]), .I1(n22));
    AND3 i2879 (.O(n3206), .I0(n780), .I1(n2789), .I2(n34));
    OR2 i2942 (.O(n3269), .I0(n3268), .I1(n3267));
    AND3 i2944 (.O(n3271), .I0(n32_adj_32), .I1(led_row_c_1), .I2(n39));
    OR2 i2945 (.O(n3272), .I0(n3271), .I1(n3270));
    OR2 i1_adj_21 (.O(n78_adj_7), .I0(n70_adj_9), .I1(n67_adj_8));
    AND2 i1_adj_22 (.O(col3[3]), .I0(n792), .I1(n23));
    AND2 i2947 (.O(n3274), .I0(scan_data[2]), .I1(n27_adj_27));
    OR2 i1_adj_23 (.O(n81_adj_10), .I0(n76_adj_6), .I1(n73_adj_3));
    OR2 i2948 (.O(n3275), .I0(n3274), .I1(n3273));
    AND6 i2883 (.O(n3210), .I0(n4_adj_67), .I1(scan_data[3]), .I2(n832), 
         .I3(n5_adj_69), .I4(led_row_c_5), .I5(n15));
    AND3 i2950 (.O(n3277), .I0(n3293), .I1(led_row_c_3), .I2(n37));
    OR2 i2951 (.O(n3278), .I0(n3277), .I1(n3276));
    OR2 i2884 (.O(n3211), .I0(n3210), .I1(n3209));
    AND2 i2953 (.O(n3280), .I0(scan_data[3]), .I1(scan_data[2]));
    AND5 i2886 (.O(n3213), .I0(n10_adj_70), .I1(n14_adj_41), .I2(n832), 
         .I3(led_row_c_6), .I4(n2784));
    OR2 i2954 (.O(n20), .I0(n3280), .I1(n3279));
    OR2 i2887 (.O(n3214), .I0(n3213), .I1(n3212));
    AND2 i2956 (.O(n3283), .I0(scan_data[2]), .I1(n6_adj_28));
    AND4 i2889 (.O(n3216), .I0(n11), .I1(n6_adj_74), .I2(n3215), .I3(led_row_c_2));
    OR2 i2957 (.O(n3284), .I0(n3283), .I1(n3282));
    AND2 i2959 (.O(n3286), .I0(scan_data[0]), .I1(n28_adj_47));
    AND2 i2890 (.O(n3217), .I0(led_row_c_3), .I1(n32));
    OR2 i2960 (.O(n3287), .I0(n3286), .I1(n3285));
    OR2 i2891 (.O(n3218), .I0(n3217), .I1(n3216));
    AND3 i2893 (.O(n3220), .I0(n4_adj_76), .I1(led_row_c_1), .I2(n32_adj_29));
    AND2 i2367 (.O(n2698), .I0(n2691), .I1(cnt_next[18]));
    AND2 i2085 (.O(n2416), .I0(n2407), .I1(scan_data[1]));
    AND2 i2962 (.O(n3289), .I0(scan_data[3]), .I1(n4_adj_67));
    OR2 i2963 (.O(n3290), .I0(n3289), .I1(n3288));
    AND2 i2965 (.O(n3292), .I0(scan_data[3]), .I1(n22));
    OR2 i2966 (.O(n3293), .I0(n3292), .I1(n3291));
    AND2 i2968 (.O(n3295), .I0(scan_data[1]), .I1(n21_adj_49));
    OR2 i2969 (.O(n3296), .I0(n3295), .I1(n3294));
    AND2 i2971 (.O(n3298), .I0(scan_data[2]), .I1(n25));
    OR2 i2972 (.O(n3299), .I0(n3298), .I1(n3297));
    AND2 i2974 (.O(n3301), .I0(scan_data[3]), .I1(n4_adj_67));
    OR2 i2975 (.O(n3302), .I0(n3301), .I1(n3300));
    AND2 i2977 (.O(n3304), .I0(scan_data[2]), .I1(n6_adj_28));
    OR2 i2978 (.O(n3305), .I0(n3304), .I1(n3303));
    AND2 i2980 (.O(n3307), .I0(scan_data[2]), .I1(scan_data[0]));
    AND2 i2374 (.O(n2705), .I0(n2698), .I1(cnt_next[19]));
    DFFCR row_buf_i0_i7 (.Q(led_row_c_6), .D(led_row_c_5), .CLK(clk_50m_c), 
          .CE(n847), .R(reset_n_c));   // led.v(26[13] 35[11])
    DFFCR row_buf_i0_i6 (.Q(led_row_c_5), .D(led_row_c_4), .CLK(clk_50m_c), 
          .CE(n847), .R(reset_n_c));   // led.v(26[13] 35[11])
    DFFCR row_buf_i0_i5 (.Q(led_row_c_4), .D(led_row_c_3), .CLK(clk_50m_c), 
          .CE(n847), .R(reset_n_c));   // led.v(26[13] 35[11])
    DFFCR row_buf_i0_i4 (.Q(led_row_c_3), .D(led_row_c_2), .CLK(clk_50m_c), 
          .CE(n847), .R(reset_n_c));   // led.v(26[13] 35[11])
    DFFCR row_buf_i0_i3 (.Q(led_row_c_2), .D(led_row_c_1), .CLK(clk_50m_c), 
          .CE(n847), .R(reset_n_c));   // led.v(26[13] 35[11])
    DFFCR row_buf_i0_i2 (.Q(led_row_c_1), .D(led_row_c_0), .CLK(clk_50m_c), 
          .CE(n847), .R(reset_n_c));   // led.v(26[13] 35[11])
    DFFR cnt_next_152_153__i25 (.Q(cnt_next[24]), .D(n133), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    AND2 i1_adj_24 (.O(n3152), .I0(n3150), .I1(n3362));
    OR2 i2981 (.O(n3308), .I0(n3307), .I1(n3306));
    DFFR cnt_next_152_153__i24 (.Q(cnt_next[23]), .D(n134), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i23 (.Q(cnt_next[22]), .D(n135), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i22 (.Q(cnt_next[21]), .D(n136), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i21 (.Q(cnt_next[20]), .D(n137), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i20 (.Q(cnt_next[19]), .D(n138), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i19 (.Q(cnt_next[18]), .D(n139), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i18 (.Q(cnt_next[17]), .D(n140), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i17 (.Q(cnt_next[16]), .D(n141), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i16 (.Q(cnt_next[15]), .D(n142), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i15 (.Q(cnt_next[14]), .D(n143), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i14 (.Q(cnt_next[13]), .D(n144), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i13 (.Q(cnt_next[12]), .D(n145), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i12 (.Q(cnt_next[11]), .D(n146), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i11 (.Q(cnt_next[10]), .D(n147), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i10 (.Q(cnt_next[9]), .D(n148), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i9 (.Q(cnt_next[8]), .D(n149), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i8 (.Q(cnt_next[7]), .D(n150), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i7 (.Q(cnt_next[6]), .D(n151), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i6 (.Q(cnt_next[5]), .D(n152), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i5 (.Q(cnt_next[4]), .D(n153), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i4 (.Q(cnt_next[3]), .D(n154), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i3 (.Q(cnt_next[2]), .D(n155), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_next_152_153__i2 (.Q(cnt_next[1]), .D(n156), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    DFFR cnt_scan_155__i15 (.Q(cnt_scan[15]), .D(n70_adj_68), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(28[23:33])
    DFFR cnt_scan_155__i14 (.Q(cnt_scan[14]), .D(n71), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(28[23:33])
    DFFR scan_data_154__i0 (.Q(scan_data[0]), .D(n2778), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(53[24:38])
    DFFR cnt_scan_155__i13 (.Q(cnt_scan[13]), .D(n72), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(28[23:33])
    DFFR cnt_scan_155__i12 (.Q(cnt_scan[12]), .D(n73_adj_79), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(28[23:33])
    DFFR cnt_scan_155__i11 (.Q(cnt_scan[11]), .D(n74), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(28[23:33])
    DFFR cnt_scan_155__i10 (.Q(cnt_scan[10]), .D(n75), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(28[23:33])
    DFFR cnt_scan_155__i9 (.Q(cnt_scan[9]), .D(n76_adj_80), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(28[23:33])
    DFFR cnt_scan_155__i8 (.Q(cnt_scan[8]), .D(n77), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(28[23:33])
    DFFR cnt_scan_155__i7 (.Q(cnt_scan[7]), .D(n78_adj_55), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(28[23:33])
    DFFR cnt_scan_155__i6 (.Q(cnt_scan[6]), .D(n79), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(28[23:33])
    DFFR cnt_scan_155__i5 (.Q(cnt_scan[5]), .D(n80), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(28[23:33])
    DFFR cnt_scan_155__i4 (.Q(cnt_scan[4]), .D(n81_adj_64), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(28[23:33])
    DFFR cnt_scan_155__i3 (.Q(cnt_scan[3]), .D(n82), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(28[23:33])
    DFFR cnt_scan_155__i2 (.Q(cnt_scan[2]), .D(n83), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(28[23:33])
    IBUF reset_n_pad (.O(reset_n_c), .I0(reset_n));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(186[8:12])
    INV i2888 (.O(n3215), .I0(led_row_c_3));
    AND2 i2177 (.O(n2508), .I0(n2501), .I1(cnt_scan[7]));
    AND4 i2870 (.O(n3197), .I0(led_row_c_4), .I1(n805), .I2(n2784), 
         .I3(n3299));
    AND2 i1_adj_25 (.O(n3153), .I0(n3150), .I1(n3338));
    OR2 i2828 (.O(n3157), .I0(n1685), .I1(led_row_c_4));
    AND2 i2983 (.O(n3310), .I0(scan_data[2]), .I1(n4));
    AND2 i2381 (.O(n2712), .I0(n2705), .I1(cnt_next[20]));
    AND2 i2_adj_26 (.O(n76_adj_6), .I0(n7_adj_66), .I1(n3202));
    AND2 i2_adj_27 (.O(n73_adj_3), .I0(n4_adj_54), .I1(n3199));
    DFFR cnt_scan_155__i1 (.Q(cnt_scan[1]), .D(n84), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(28[23:33])
    INV i1252 (.O(n7_adj_65), .I0(n1588));
    DFFR scan_data_154__i6 (.Q(scan_data[6]), .D(n34_adj_63), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(53[24:38])
    INV i1349 (.O(n805), .I0(n1685));
    DFFR scan_data_154__i5 (.Q(scan_data[5]), .D(n35), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(53[24:38])
    DFFR scan_data_154__i4 (.Q(scan_data[4]), .D(n36), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(53[24:38])
    DFFR scan_data_154__i3 (.Q(scan_data[3]), .D(n37_adj_62), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(53[24:38])
    DFFR scan_data_154__i2 (.Q(scan_data[2]), .D(n38), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(53[24:38])
    DFFR scan_data_154__i1 (.Q(scan_data[1]), .D(n39_adj_60), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(53[24:38])
    DFFR cnt_next_152_153__i1 (.Q(cnt_next[0]), .D(n157), .CLK(clk_50m_c), 
         .R(reset_n_c)) /* synthesis syn_use_carry_chain=1 */ ;   // led.v(48[23:33])
    OR2 i2984 (.O(n3311), .I0(n3310), .I1(n3309));
    AND2 i2388 (.O(n2719), .I0(n2712), .I1(cnt_next[21]));
    DFFCR row_buf_i0_i1 (.Q(led_row_c_0), .D(led_row_c_7), .CLK(clk_50m_c), 
          .CE(n847), .R(reset_n_c));   // led.v(26[13] 35[11])
    OBUF led_col_pad_7 (.O(led_col[7]), .I0(col_buf[7]));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    AND2 i2106 (.O(n2437), .I0(n2430), .I1(scan_data[4]));
    AND2 i2986 (.O(n3313), .I0(scan_data[0]), .I1(n28_adj_47));
    IBUF clk_50m_pad (.O(clk_50m_c), .I0(clk_50m));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(186[8:12])
    OBUF led_row_pad_0 (.O(led_row[0]), .I0(led_row_c_0));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    AND2 i2_adj_28 (.O(n70_adj_9), .I0(n7_adj_65), .I1(n3218));
    OBUF led_row_pad_1 (.O(led_row[1]), .I0(led_row_c_1));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF led_row_pad_2 (.O(led_row[2]), .I0(led_row_c_2));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OR2 i2987 (.O(n3314), .I0(n3313), .I1(n3312));
    AND3 i2989 (.O(n3316), .I0(n18_adj_53), .I1(scan_data[0]), .I2(n4));
    OBUF led_row_pad_3 (.O(led_row[3]), .I0(led_row_c_3));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF led_row_pad_4 (.O(led_row[4]), .I0(led_row_c_4));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF led_row_pad_5 (.O(led_row[5]), .I0(led_row_c_5));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OR2 i2990 (.O(n3317), .I0(n3316), .I1(n3315));
    AND2 i2992 (.O(n3319), .I0(scan_data[3]), .I1(n7));
    INV i2467 (.O(n4_adj_67), .I0(n18_adj_53));
    AND2 i1341 (.O(n157), .I0(n49), .I1(n130));
    INV i1236 (.O(n8_adj_72), .I0(n1572));
    OBUF led_row_pad_6 (.O(led_row[6]), .I0(led_row_c_6));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF led_row_pad_7 (.O(led_row[7]), .I0(led_row_c_7));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF led_col_pad_0 (.O(led_col[0]), .I0(col_buf[0]));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    AND2 i2283 (.O(n2614), .I0(n2607), .I1(cnt_next[6]));
    OR2 i2993 (.O(n3320), .I0(n3319), .I1(n3318));
    OBUF led_col_pad_1 (.O(led_col[1]), .I0(col_buf[1]));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF led_col_pad_2 (.O(led_col[2]), .I0(col_buf[2]));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF led_col_pad_3 (.O(led_col[3]), .I0(col_buf[3]));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    AND2 i2995 (.O(n3322), .I0(scan_data[3]), .I1(n12));
    OR2 i2838 (.O(n3167), .I0(n1719), .I1(led_row_c_4));
    AND2 i2_adj_29 (.O(n67_adj_8), .I0(n8), .I1(n3221));
    OBUF led_col_pad_4 (.O(led_col[4]), .I0(col_buf[4]));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    AND2 i2113 (.O(n2444), .I0(n2437), .I1(scan_data[5]));
    AND2 i2092 (.O(n2423), .I0(n2416), .I1(scan_data[2]));
    OR2 i2894 (.O(n3221), .I0(n3220), .I1(n3219));
    OBUF led_col_pad_5 (.O(led_col[5]), .I0(col_buf[5]));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF led_col_pad_6 (.O(led_col[6]), .I0(col_buf[6]));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    XOR2 i2082 (.O(n39_adj_60), .I0(n2407), .I1(scan_data[1]));
    AND2 i2876 (.O(n3203), .I0(n14), .I1(n8_adj_16));
    AND2 i2395 (.O(n2726), .I0(n2719), .I1(cnt_next[22]));
    AND2 i2402 (.O(n2733), .I0(n2726), .I1(cnt_next[23]));
    AND2 i2304 (.O(n2635), .I0(n2628), .I1(cnt_next[9]));
    AND2 i2269 (.O(n2600), .I0(n2593), .I1(cnt_next[4]));
    XOR2 i2089 (.O(n38), .I0(n2416), .I1(scan_data[2]));
    XOR2 i2139 (.O(n83), .I0(n2466), .I1(cnt_scan[2]));
    OR2 i2996 (.O(n3323), .I0(n3322), .I1(n3321));
    AND2 i2998 (.O(n3325), .I0(scan_data[3]), .I1(n18_adj_44));
    OR2 i2999 (.O(n3326), .I0(n3325), .I1(n3324));
    AND2 i3001 (.O(n3328), .I0(scan_data[0]), .I1(scan_data[1]));
    XOR2 i2252 (.O(n128), .I0(n2579), .I1(cnt_next[2]));
    OR2 i1_adj_30 (.O(n12_adj_71), .I0(n1695), .I1(scan_data[3]));
    OR2 i3002 (.O(n3329), .I0(n3328), .I1(n3327));
    AND2 i3004 (.O(n3331), .I0(scan_data[1]), .I1(n22));
    OR2 i3005 (.O(n3332), .I0(n3331), .I1(n3330));
    AND3 i3007 (.O(n3334), .I0(n3314), .I1(led_row_c_5), .I2(n28));
    OR2 i3008 (.O(n3335), .I0(n3334), .I1(n3333));
    OR2 i1_adj_31 (.O(n3156), .I0(n1695), .I1(scan_data[1]));
    AND2 i2149 (.O(n2480), .I0(n2473), .I1(cnt_scan[3]));
    AND3 i3010 (.O(n3337), .I0(n30), .I1(led_row_c_1), .I2(n39));
    OR2 i3011 (.O(n3338), .I0(n3337), .I1(n3336));
    AND3 i3013 (.O(n3340), .I0(n3359), .I1(led_row_c_7), .I2(n10));
    OR2 i3014 (.O(n3341), .I0(n3340), .I1(n3339));
    AND2 i2262 (.O(n2593), .I0(n2586), .I1(cnt_next[3]));
    XOR2 i2096 (.O(n37_adj_62), .I0(n2423), .I1(scan_data[3]));
    AND2 i3016 (.O(n3343), .I0(scan_data[0]), .I1(scan_data[1]));
    AND2 i2248 (.O(n2579), .I0(cnt_next[0]), .I1(cnt_next[1]));
    XOR2 i2103 (.O(n36), .I0(n2430), .I1(scan_data[4]));
    OR2 i1344 (.O(n1681), .I0(n18_adj_53), .I1(scan_data[0]));
    AND2 i2255 (.O(n2586), .I0(n2579), .I1(cnt_next[2]));
    AND2 i3019 (.O(n3346), .I0(scan_data[3]), .I1(n18_adj_44));
    OR2 i1348 (.O(n1685), .I0(n1572), .I1(n1606));
    AND2 i2135 (.O(n2466), .I0(cnt_scan[0]), .I1(cnt_scan[1]));
    INV i1250 (.O(n4_adj_54), .I0(n1586));
    INV i2829 (.O(n5_adj_86), .I0(n3157));
    AND2 i2290 (.O(n2621), .I0(n2614), .I1(cnt_next[7]));
    OR2 i3020 (.O(n3347), .I0(n3346), .I1(n3345));
    XOR2 i2245 (.O(n129), .I0(cnt_next[0]), .I1(cnt_next[1]));
    INV i1246 (.O(n7_adj_66), .I0(n1582));
    INV i1244 (.O(n8), .I0(n1580));
    AND2 i2142 (.O(n2473), .I0(n2466), .I1(cnt_scan[2]));
    AND2 i3022 (.O(n3349), .I0(scan_data[2]), .I1(n6_adj_50));
    XOR2 i2132 (.O(n84), .I0(cnt_scan[0]), .I1(cnt_scan[1]));
    OR2 i3023 (.O(n3350), .I0(n3349), .I1(n3348));
    XOR2 i2110 (.O(n35), .I0(n2437), .I1(scan_data[5]));
    OR2 i1358 (.O(n1695), .I0(scan_data[4]), .I1(n1606));
    AND2 i2871 (.O(n3198), .I0(led_row_c_5), .I1(n48));
    OR2 i1362 (.O(n1699), .I0(n1685), .I1(led_row_c_0));
    XOR2 i2266 (.O(n126), .I0(n2593), .I1(cnt_next[4]));
    XOR2 i2273 (.O(n125), .I0(n2600), .I1(cnt_next[5]));
    AND4 i3025 (.O(n3352), .I0(n10), .I1(n3356), .I2(led_row_c_7), .I3(n15));
    OR2 i1249 (.O(n1586), .I0(led_row_c_6), .I1(led_row_c_7));
    OR2 i1239 (.O(n1576), .I0(n846), .I1(led_row_c_4));
    OR2 i3026 (.O(n3353), .I0(n3352), .I1(n3351));
    XOR2 i2280 (.O(n124), .I0(n2607), .I1(cnt_next[6]));
    AND3 i3028 (.O(n3355), .I0(n1628), .I1(scan_data[2]), .I2(n4));
    XOR2 i2153 (.O(n81_adj_64), .I0(n2480), .I1(cnt_scan[4]));
    OR2 i3029 (.O(n3356), .I0(n3355), .I1(n3354));
    XOR2 i2160 (.O(n80), .I0(n2487), .I1(cnt_scan[5]));
    AND2 i3031 (.O(n3358), .I0(scan_data[3]), .I1(n4_adj_67));
    OR2 i3032 (.O(n3359), .I0(n3358), .I1(n3357));
    AND2 i1372 (.O(n1709), .I0(n1656), .I1(n1681));
    XOR2 i2117 (.O(n34_adj_63), .I0(n2444), .I1(scan_data[6]));
    AND2 i2184 (.O(n2515), .I0(n2508), .I1(cnt_scan[8]));
    XOR2 i2287 (.O(n123), .I0(n2614), .I1(cnt_next[7]));
    XOR2 i2294 (.O(n122), .I0(n2621), .I1(cnt_next[8]));
    OR2 i1380 (.O(n1717), .I0(n1695), .I1(led_row_c_2));
    AND3 i3034 (.O(n3361), .I0(n30_adj_40), .I1(led_row_c_1), .I2(n39));
    XOR2 i2167 (.O(n79), .I0(n2494), .I1(cnt_scan[6]));
    AND2 i2170 (.O(n2501), .I0(n2494), .I1(cnt_scan[6]));
    XOR2 i2174 (.O(n78_adj_55), .I0(n2501), .I1(cnt_scan[7]));
    XOR2 i2301 (.O(n121), .I0(n2628), .I1(cnt_next[9]));
    XOR2 i2308 (.O(n120), .I0(n2635), .I1(cnt_next[10]));
    OR2 i3035 (.O(n3362), .I0(n3361), .I1(n3360));
    AND3 i3037 (.O(n3364), .I0(n19), .I1(scan_data[3]), .I2(n22));
    OR2 i3038 (.O(n3365), .I0(n3364), .I1(n3363));
    XOR2 i2181 (.O(n77), .I0(n2508), .I1(cnt_scan[8]));
    XOR2 i2315 (.O(n119), .I0(n2642), .I1(cnt_next[11]));
    XOR2 i2188 (.O(n76_adj_80), .I0(n2515), .I1(cnt_scan[9]));
    OR2 i1_adj_32 (.O(n846), .I0(n844), .I1(n8_adj_73));
    AND2 i1_adj_33 (.O(n816), .I0(n812), .I1(n81_adj_2));
    AND2 i1_adj_34 (.O(n836), .I0(n835), .I1(n6_adj_28));
    AND2 i1_adj_35 (.O(n835), .I0(n31), .I1(scan_data[0]));
    XOR2 i2259 (.O(n127), .I0(n2586), .I1(cnt_next[3]));
    OR6 i1_adj_36 (.O(n49), .I0(n14_adj_90), .I1(cnt_next[10]), .I2(n12_adj_97), 
        .I3(n13), .I4(n776), .I5(cnt_next[20]));
    AND2 i1_adj_37 (.O(n817), .I0(n812), .I1(n81_adj_13));
    AND2 i2163 (.O(n2494), .I0(n2487), .I1(cnt_scan[5]));
    XOR2 i2322 (.O(n118), .I0(n2649), .I1(cnt_next[12]));
    AND2 i1_adj_38 (.O(n818), .I0(n812), .I1(n81));
    OR2 i1277 (.O(n1614), .I0(scan_data[0]), .I1(scan_data[2]));
    XOR2 i2329 (.O(n117), .I0(n2656), .I1(cnt_next[13]));
    XOR2 i2195 (.O(n75), .I0(n2522), .I1(cnt_scan[10]));
    OR2 i1342 (.O(n1679), .I0(n1582), .I1(n1586));
    OR2 scan_data_6__I_0_67_i8 (.O(n8_adj_73), .I0(scan_data[2]), .I1(n6_adj_28));
    AND2 i1_adj_39 (.O(n785), .I0(n784), .I1(n78_adj_7));
    AND2 i1_adj_40 (.O(n786), .I0(n784), .I1(n78_adj_12));
    AND2 i1_adj_41 (.O(n819), .I0(n812), .I1(n81_adj_10));
    OR2 scan_data_6__I_0_67_i11 (.O(n1606), .I0(scan_data[6]), .I1(scan_data[5]));
    AND3 i2_adj_42 (.O(n2764), .I0(n4_adj_54), .I1(n3248), .I2(n805));
    AND2 i3036 (.O(n3363), .I0(n4), .I1(n12_adj_95));
    AND2 i5 (.O(col4[7]), .I0(n805), .I1(n5));
    XOR2 i2146 (.O(n82), .I0(n2473), .I1(cnt_scan[3]));
    OR2 i1382 (.O(n1719), .I0(n1695), .I1(scan_data[2]));
    AND3 i3033 (.O(n3360), .I0(n3317), .I1(n14), .I2(led_row_c_0));
    AND2 i1_adj_43 (.O(n5), .I0(scan_data[0]), .I1(scan_data[2]));
    AND2 i3030 (.O(n3357), .I0(n4), .I1(n5));
    AND2 i1_adj_44 (.O(n787), .I0(n784), .I1(n78_adj_4));
    AND3 i3027 (.O(n3354), .I0(n19), .I1(n22), .I2(scan_data[3]));
    XOR2 i28 (.O(n31), .I0(scan_data[3]), .I1(scan_data[2]));
    AND4 i3024 (.O(n3351), .I0(n8_adj_72), .I1(n20_adj_59), .I2(n2789), 
         .I3(led_row_c_6));
    AND2 i3021 (.O(n3348), .I0(n22), .I1(n25));
    AND2 i2_adj_45 (.O(n2757), .I0(n4_adj_81), .I1(n3353));
    AND2 i3018 (.O(n3345), .I0(n4), .I1(n3350));
    AND2 i3015 (.O(n3342), .I0(n11), .I1(scan_data[2]));
    AND3 i3012 (.O(n3339), .I0(n25_adj_61), .I1(n2789), .I2(led_row_c_6));
    AND3 i3009 (.O(n3336), .I0(n3320), .I1(n14), .I2(led_row_c_0));
    AND2 i2_adj_46 (.O(n76_adj_11), .I0(n7_adj_66), .I1(n3208));
    AND3 i3006 (.O(n3333), .I0(n3365), .I1(n2784), .I2(led_row_c_4));
    OR2 i1_adj_47 (.O(n20_adj_59), .I0(n14_adj_43), .I1(n22));
    AND2 i3003 (.O(n3330), .I0(n6_adj_28), .I1(n23_adj_58));
    AND2 i3000 (.O(n3327), .I0(n11), .I1(n22));
    OR2 i1_adj_48 (.O(n23_adj_58), .I0(n11), .I1(scan_data[2]));
    OR2 i1_adj_49 (.O(n34), .I0(n836), .I1(n726));
    AND2 i2_adj_50 (.O(n67), .I0(n8), .I1(n3205));
    OR3 i2_adj_51 (.O(n845), .I0(scan_data[1]), .I1(n844), .I2(n22));
    AND2 i2997 (.O(n3324), .I0(n4), .I1(n3329));
    AND2 i1_adj_52 (.O(n824), .I0(n805), .I1(scan_data[2]));
    AND2 i12 (.O(n28_adj_98), .I0(n24), .I1(n23_adj_46));
    AND2 i2994 (.O(n3321), .I0(n4), .I1(n5));
    AND2 i2991 (.O(n3318), .I0(n4), .I1(n5));
    OR3 i1319 (.O(n1656), .I0(n3343), .I1(n3342), .I2(scan_data[3]));
    INV i2843 (.O(n3150), .I0(n3171));
    AND2 i1318 (.O(n156), .I0(n49), .I1(n129));
    AND2 i1317 (.O(n155), .I0(n49), .I1(n128));
    AND2 i1316 (.O(n154), .I0(n49), .I1(n127));
    INV i2848 (.O(n3175), .I0(n786));
    AND2 i1315 (.O(n153), .I0(n49), .I1(n126));
    INV i2849 (.O(n3176), .I0(n813));
    INV i2851 (.O(n3178), .I0(n785));
    INV i2852 (.O(n3179), .I0(n819));
    AND2 i2_adj_53 (.O(n70_adj_1), .I0(n7_adj_65), .I1(n3230));
    OR2 i1_adj_54 (.O(n18_adj_53), .I0(scan_data[1]), .I1(scan_data[2]));
    AND2 i1314 (.O(n152), .I0(n49), .I1(n125));
    INV i2854 (.O(n3181), .I0(n788));
    AND2 i1313 (.O(n151), .I0(n49), .I1(n124));
    INV i2855 (.O(n3182), .I0(n816));
    AND2 i1312 (.O(n150), .I0(n49), .I1(n123));
    AND2 i1311 (.O(n149), .I0(n49), .I1(n122));
    AND2 i2_adj_55 (.O(n73), .I0(n4_adj_54), .I1(n3227));
    INV i2857 (.O(n3184), .I0(n787));
    AND2 i1310 (.O(n148), .I0(n49), .I1(n121));
    AND2 i1309 (.O(n147), .I0(n49), .I1(n120));
    AND2 i1308 (.O(n146), .I0(n49), .I1(n119));
    INV i2858 (.O(n3185), .I0(n818));
    AND2 i1307 (.O(n145), .I0(n49), .I1(n118));
    INV i2860 (.O(n3187), .I0(n791));
    AND2 i1306 (.O(n144), .I0(n49), .I1(n117));
    AND2 i1305 (.O(n143), .I0(n49), .I1(n116));
    AND2 i2_adj_56 (.O(n76), .I0(n7_adj_66), .I1(n3224));
    INV i2861 (.O(n3188), .I0(n817));
    AND2 i1304 (.O(n142), .I0(n49), .I1(n115));
    AND2 i1303 (.O(n141), .I0(n49), .I1(n114));
    OR2 i1_adj_57 (.O(n15_adj_51), .I0(n11), .I1(scan_data[3]));
    AND2 i1302 (.O(n140), .I0(n49), .I1(n113));
    AND2 i1301 (.O(n139), .I0(n49), .I1(n112));
    AND2 i1300 (.O(n138), .I0(n49), .I1(n111));
    AND2 i1299 (.O(n137), .I0(n49), .I1(n110));
    AND2 i1298 (.O(n136), .I0(n49), .I1(n109));
    AND2 i1297 (.O(n135), .I0(n49), .I1(n108));
    AND2 i1296 (.O(n134), .I0(n49), .I1(n107));
    AND3 i2988 (.O(n3315), .I0(n22), .I1(n11), .I2(scan_data[3]));
    INV i2863 (.O(n3190), .I0(n790));
    INV i2864 (.O(n3191), .I0(n815));
    INV i2866 (.O(n3193), .I0(n789));
    AND3 i2985 (.O(n3312), .I0(n31), .I1(n11), .I2(scan_data[1]));
    AND2 i2982 (.O(n3309), .I0(n22), .I1(scan_data[0]));
    XOR2 i324 (.O(n659), .I0(led_row_c_3), .I1(led_row_c_2));
    INV i2867 (.O(n3194), .I0(n814));
    AND6 i15_adj_58 (.O(n2748), .I0(n28_adj_82), .I1(cnt_next[19]), .I2(n18_adj_93), 
         .I3(n26_adj_84), .I4(n27_adj_83), .I5(cnt_next[0]));
    AND2 i2979 (.O(n3306), .I0(n22), .I1(n19));
    AND2 i2976 (.O(n3303), .I0(n22), .I1(n6_adj_50));
    INV i2869 (.O(n3196), .I0(n49));
    AND2 i2198 (.O(n2529), .I0(n2522), .I1(cnt_scan[10]));
    AND2 i2_adj_59 (.O(n18_adj_93), .I0(cnt_next[3]), .I1(cnt_next[15]));
    XOR2 i2336 (.O(n116), .I0(n2663), .I1(cnt_next[14]));
    AND2 i3 (.O(n19_adj_92), .I0(cnt_next[5]), .I1(cnt_next[6]));
    AND2 i4 (.O(n20_adj_91), .I0(cnt_next[16]), .I1(cnt_next[14]));
    AND2 i5_adj_60 (.O(n21_adj_89), .I0(cnt_next[9]), .I1(cnt_next[4]));
    AND2 i6 (.O(n22_adj_88), .I0(cnt_next[22]), .I1(cnt_next[1]));
    AND2 i2191 (.O(n2522), .I0(n2515), .I1(cnt_scan[9]));
    AND2 i1_adj_61 (.O(n828), .I0(n659), .I1(n7_adj_65));
    AND2 i1_adj_62 (.O(n829), .I0(n828), .I1(col4[7]));
    AND2 i2156 (.O(n2487), .I0(n2480), .I1(cnt_scan[4]));
    XOR2 i2343 (.O(n115), .I0(n2670), .I1(cnt_next[15]));
    AND3 i2_adj_63 (.O(n2760), .I0(col4[7]), .I1(n661), .I2(n4_adj_54));
    GND i2844 (.X(gnd));
    XOR2 i2202 (.O(n74), .I0(n2529), .I1(cnt_scan[11]));
    AND2 i7_adj_64 (.O(n23_adj_87), .I0(cnt_next[8]), .I1(cnt_next[23]));
    XOR2 i2350 (.O(n114), .I0(n2677), .I1(cnt_next[16]));
    XOR2 i2357 (.O(n113), .I0(n2684), .I1(cnt_next[17]));
    AND2 i8_adj_65 (.O(n24_adj_85), .I0(cnt_next[24]), .I1(cnt_next[2]));
    XOR2 i2364 (.O(n112), .I0(n2691), .I1(cnt_next[18]));
    OR2 i1281 (.O(n1618), .I0(n1588), .I1(n1580));
    AND2 i10_adj_66 (.O(n26_adj_84), .I0(n20_adj_91), .I1(n19_adj_92));
    AND2 i11_adj_67 (.O(n27_adj_83), .I0(n22_adj_88), .I1(n21_adj_89));
    AND2 i2_adj_68 (.O(n70), .I0(n7_adj_65), .I1(n3233));
    AND2 i2973 (.O(n3300), .I0(n4), .I1(n3305));
    XOR2 i2371 (.O(n111), .I0(n2698), .I1(cnt_next[19]));
    AND2 i2970 (.O(n3297), .I0(n22), .I1(n6_adj_50));
    AND2 i12_adj_69 (.O(n28_adj_82), .I0(n24_adj_85), .I1(n23_adj_87));
    INV i2243 (.O(n130), .I0(cnt_next[0]));
    INV i2130 (.O(n85), .I0(cnt_scan[0]));
    INV i2455 (.O(n2784), .I0(led_row_c_5));
    XOR2 i2378 (.O(n110), .I0(n2705), .I1(cnt_next[20]));
    OR2 i1_adj_70 (.O(n21_adj_49), .I0(scan_data[0]), .I1(n22));
    INV i1391 (.O(n775), .I0(n1727));
    XOR2 i2385 (.O(n109), .I0(n2712), .I1(cnt_next[21]));
    INV i1345 (.O(n12), .I0(n1681));
    INV scan_data_6__I_0_66_i14 (.O(col1_7__N_71), .I0(n2773));
    INV i279 (.O(n6_adj_28), .I0(scan_data[1]));
    AND2 i2967 (.O(n3294), .I0(n6_adj_28), .I1(scan_data[2]));
    XOR2 i2209 (.O(n73_adj_79), .I0(n2536), .I1(cnt_scan[12]));
    OR2 i1_adj_71 (.O(n10_adj_26), .I0(cnt_next[11]), .I1(cnt_next[21]));
    XOR2 i2392 (.O(n108), .I0(n2719), .I1(cnt_next[22]));
    XOR2 i2216 (.O(n72), .I0(n2543), .I1(cnt_scan[13]));
    INV i1343 (.O(n784), .I0(n1679));
    XOR2 i56 (.O(n27_adj_48), .I0(scan_data[2]), .I1(scan_data[1]));
    AND3 i2964 (.O(n3291), .I0(n11), .I1(n4), .I2(scan_data[2]));
    AND3 i2961 (.O(n3288), .I0(scan_data[1]), .I1(n4), .I2(scan_data[2]));
    XOR2 i2399 (.O(n107), .I0(n2726), .I1(cnt_next[23]));
    AND2 i1_adj_72 (.O(n28_adj_47), .I0(n27_adj_48), .I1(n4));
    AND2 i2205 (.O(n2536), .I0(n2529), .I1(cnt_scan[11]));
    INV scan_data_6__I_0_67_i14 (.O(col1_7__N_72), .I0(n846));
    XOR2 i2406 (.O(n106), .I0(n2733), .I1(cnt_next[24]));
    AND3 i2_adj_73 (.O(n2752), .I0(n7_adj_66), .I1(n3341), .I2(n792));
    OR2 i1390 (.O(n1727), .I0(n1624), .I1(n1717));
    INV i2839 (.O(n5_adj_56), .I0(n3167));
    AND2 i1283 (.O(n6_adj_50), .I0(scan_data[0]), .I1(scan_data[1]));
    AND3 i2_adj_74 (.O(n2770), .I0(n3275), .I1(n828), .I2(n805));
    INV i9 (.O(n22), .I0(scan_data[2]));
    AND2 i2958 (.O(n3285), .I0(n11), .I1(n3290));
    OR2 i1_adj_75 (.O(n23), .I0(n21), .I1(n18_adj_44));
    INV i3_adj_76 (.O(n15), .I0(scan_data[4]));
    INV i15_adj_77 (.O(n11), .I0(scan_data[0]));
    INV scan_data_6__I_0_69_i14 (.O(col1_7__N_74), .I0(n845));
    AND2 i1_adj_78 (.O(n831), .I0(n828), .I1(col1_7__N_71));
    INV i277 (.O(n4), .I0(scan_data[3]));
    INV i1326 (.O(n820), .I0(n3156));
    AND3 i2_adj_79 (.O(n2758), .I0(n4_adj_54), .I1(n3335), .I2(n792));
    AND2 i1_adj_80 (.O(n21), .I0(n3284), .I1(n4));
    AND2 i2_adj_81 (.O(n73_adj_15), .I0(n4_adj_54), .I1(n3236));
    INV i1373 (.O(n25_adj_61), .I0(n1709));
    AND2 i2955 (.O(n3282), .I0(n22), .I1(scan_data[0]));
    INV i1395 (.O(n776), .I0(n2748));
    AND2 i1_adj_82 (.O(n813), .I0(n812), .I1(n81_adj_5));
    OR2 i3_adj_83 (.O(n12_adj_97), .I0(cnt_next[17]), .I1(cnt_next[12]));
    AND2 i2952 (.O(n3279), .I0(n4), .I1(scan_data[1]));
    OR2 i4_adj_84 (.O(n13), .I0(cnt_next[18]), .I1(cnt_next[13]));
    INV i1292 (.O(n25), .I0(n1628));
    AND2 i2_adj_85 (.O(n18_adj_78), .I0(cnt_scan[4]), .I1(cnt_scan[1]));
    AND2 i3_adj_86 (.O(n19_adj_77), .I0(cnt_scan[13]), .I1(cnt_scan[8]));
    INV i2837 (.O(n6_adj_74), .I0(n3165));
    AND3 i2949 (.O(n3276), .I0(n31), .I1(n3215), .I2(led_row_c_2));
    AND2 i1_adj_87 (.O(n814), .I0(n812), .I1(n81_adj_22));
    OR2 i5_adj_88 (.O(n14_adj_90), .I0(n10_adj_26), .I1(cnt_next[7]));
    AND2 i1_adj_89 (.O(n780), .I0(n792), .I1(led_row_c_6));
    AND2 i4_adj_90 (.O(n20_adj_75), .I0(cnt_scan[5]), .I1(cnt_scan[3]));
    INV i1284 (.O(n14_adj_45), .I0(n6_adj_50));
    XOR2 i28_adj_91 (.O(n14_adj_43), .I0(scan_data[1]), .I1(scan_data[0]));
    AND2 i2946 (.O(n3273), .I0(n22), .I1(n19));
    OR2 i1_adj_92 (.O(n14_adj_42), .I0(scan_data[1]), .I1(n7));
    AND2 i1_adj_93 (.O(n815), .I0(n812), .I1(n81_adj_17));
    XOR2 i28_adj_94 (.O(n14_adj_41), .I0(scan_data[3]), .I1(scan_data[1]));
    AND2 i2212 (.O(n2543), .I0(n2536), .I1(cnt_scan[12]));
    AND3 i2943 (.O(n3270), .I0(n3323), .I1(n14), .I2(led_row_c_0));
    OR2 i1_adj_95 (.O(n30_adj_40), .I0(n28_adj_39), .I1(n18_adj_44));
    OR2 i1285 (.O(n1622), .I0(n20), .I1(scan_data[0]));
    AND2 i1_adj_96 (.O(n28_adj_39), .I0(n3269), .I1(n4));
    AND2 i5_adj_97 (.O(n21_adj_57), .I0(cnt_scan[12]), .I1(cnt_scan[10]));
    INV i2846 (.O(n3173), .I0(n6));
    AND2 i2940 (.O(n3267), .I0(n11), .I1(n8_adj_73));
    OR3 i1_adj_98 (.O(n30_adj_36), .I0(n3265), .I1(n3264), .I2(n28_adj_37));
    AND2 i1287 (.O(n1624), .I0(n1622), .I1(n18_adj_53));
    INV i1282 (.O(n812), .I0(n1618));
    AND2 i1_adj_99 (.O(n28_adj_37), .I0(n27_adj_38), .I1(n22));
    AND2 i1_adj_100 (.O(n832), .I0(n14), .I1(scan_data[0]));
    INV i2835 (.O(n4_adj_76), .I0(n3163));
    AND2 i2937 (.O(n3264), .I0(n6_adj_28), .I1(n5));
    OR2 i1_adj_101 (.O(n27_adj_38), .I0(n11), .I1(scan_data[1]));
    XOR2 i2223 (.O(n71), .I0(n2550), .I1(cnt_scan[14]));
    INV i2833 (.O(n4_adj_94), .I0(n3161));
    OR2 i1_adj_102 (.O(n32_adj_32), .I0(n30_adj_33), .I1(n27_adj_35));
    AND2 i1_adj_103 (.O(n30_adj_33), .I0(n29_adj_34), .I1(n22));
    OR2 i1_adj_104 (.O(n29_adj_34), .I0(n6_adj_28), .I1(n18));
    AND2 i1_adj_105 (.O(n27_adj_35), .I0(n3263), .I1(n4));
    AND2 i2_adj_106 (.O(n67_adj_18), .I0(n8), .I1(n3245));
    AND2 i2934 (.O(n3261), .I0(n22), .I1(scan_data[0]));
    AND2 i1_adj_107 (.O(n18), .I0(n11), .I1(scan_data[3]));
    OR2 i1_adj_108 (.O(n32_adj_29), .I0(n30_adj_31), .I1(n27_adj_30));
    INV equal_260_i50 (.O(n465), .I0(n49));
    OR2 i1_adj_109 (.O(n29), .I0(n6_adj_28), .I1(scan_data[3]));
    AND2 i2931 (.O(n3258), .I0(n22), .I1(scan_data[0]));
    AND2 i1_adj_110 (.O(n27_adj_30), .I0(n3260), .I1(n4));
    OR2 i1291 (.O(n1628), .I0(scan_data[0]), .I1(scan_data[1]));
    XOR2 i2230 (.O(n70_adj_68), .I0(n2557), .I1(cnt_scan[15]));
    INV i1242 (.O(n32), .I0(n1578));
    AND2 i6_adj_111 (.O(n22_adj_52), .I0(cnt_scan[7]), .I1(cnt_scan[2]));
    INV i1278 (.O(n7), .I0(n1614));
    AND3 i2873 (.O(n3200), .I0(n780), .I1(n2789), .I2(n3326));
    INV i1270 (.O(n5_adj_69), .I0(n1606));
    INV i42 (.O(n10), .I0(led_row_c_6));
    AND2 i2219 (.O(n2550), .I0(n2543), .I1(cnt_scan[13]));
    AND2 i1295 (.O(n133), .I0(n49), .I1(n106));
    AND2 i1_adj_112 (.O(n33), .I0(n3257), .I1(n4));
    OR2 i1_adj_113 (.O(n30), .I0(n33), .I1(n18_adj_44));
    AND2 i2226 (.O(n2557), .I0(n2550), .I1(cnt_scan[14]));
    AND2 i2928 (.O(n3255), .I0(n22), .I1(n27_adj_27));
    AND2 i2925 (.O(n3252), .I0(n14), .I1(n8_adj_16));
    OR2 i1_adj_114 (.O(n27_adj_27), .I0(scan_data[0]), .I1(n6_adj_28));
    XOR2 i1_adj_115 (.O(n2778), .I0(scan_data[0]), .I1(n3196));
    AND2 i1_adj_116 (.O(n8_adj_16), .I0(col1_7__N_74), .I1(led_row_c_0));
    OR2 i2872 (.O(n3199), .I0(n3198), .I1(n3197));
    OR2 i1_adj_117 (.O(n81_adj_22), .I0(n76_adj_25), .I1(n2760));
    OR2 i1_adj_118 (.O(n78_adj_24), .I0(n829), .I1(n67_adj_23));
    AND2 i2276 (.O(n2607), .I0(n2600), .I1(cnt_next[5]));
    AND2 i2_adj_119 (.O(n73_adj_21), .I0(n4_adj_54), .I1(n3242));
    AND4 i2922 (.O(n3249), .I0(led_row_c_6), .I1(n835), .I2(n2789), 
         .I3(n820));
    AND3 i2919 (.O(n3246), .I0(n3296), .I1(n2784), .I2(led_row_c_4));
    AND2 i2916 (.O(n3243), .I0(n14), .I1(n8_adj_16));
    AND3 i2913 (.O(n3240), .I0(col1_7__N_71), .I1(n2784), .I2(led_row_c_4));
    INV i39 (.O(n39), .I0(led_row_c_0));
    INV i38 (.O(n14), .I0(led_row_c_1));
    AND2 i2874 (.O(n3201), .I0(led_row_c_7), .I1(n64));
    INV i37 (.O(n37), .I0(led_row_c_2));
    INV i28_adj_120 (.O(n28), .I0(led_row_c_4));
    OR2 i1_adj_121 (.O(n81_adj_17), .I0(n76_adj_20), .I1(n73_adj_21));
    OR2 i1_adj_122 (.O(n78_adj_19), .I0(n831), .I1(n67_adj_18));
    AND2 i2_adj_123 (.O(n76_adj_20), .I0(n7_adj_66), .I1(n3239));
    AND2 i1_adj_124 (.O(n788), .I0(n784), .I1(n78));
    AND3 i2910 (.O(n3237), .I0(n780), .I1(n2789), .I2(n3347));
    AND2 i1_adj_125 (.O(n789), .I0(n784), .I1(n78_adj_24));
    
endmodule
//
// Verilog Description of module AND2
// module not written out since it is a black-box. 
//

//
// Verilog Description of module OR2
// module not written out since it is a black-box. 
//

//
// Verilog Description of module OR3
// module not written out since it is a black-box. 
//

//
// Verilog Description of module XOR2
// module not written out since it is a black-box. 
//

//
// Verilog Description of module AND4
// module not written out since it is a black-box. 
//

//
// Verilog Description of module AND3
// module not written out since it is a black-box. 
//

//
// Verilog Description of module AND6
// module not written out since it is a black-box. 
//

//
// Verilog Description of module VCC
// module not written out since it is a black-box. 
//

//
// Verilog Description of module INV
// module not written out since it is a black-box. 
//

//
// Verilog Description of module AND5
// module not written out since it is a black-box. 
//

//
// Verilog Description of module OR6
// module not written out since it is a black-box. 
//

//
// Verilog Description of module GND
// module not written out since it is a black-box. 
//

