// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Mon May 29 00:01:31 2023
//
// Verilog Description of module CALCULATE
//

module CALCULATE (clk, reset, key_in, PointTime, led_int_Data0, led_int_Data1, 
            led_int_Data2, key_out) /* synthesis syn_module_defined=1 */ ;   // calculate.v(1[8:17])
    input clk;   // calculate.v(3[11:14])
    input reset;   // calculate.v(3[15:20])
    input [3:0]key_in;   // calculate.v(4[17:23])
    output PointTime;   // calculate.v(5[12:21])
    output [3:0]led_int_Data0;   // calculate.v(6[18:31])
    output [3:0]led_int_Data1;   // calculate.v(7[18:31])
    output [3:0]led_int_Data2;   // calculate.v(8[18:31])
    output [3:0]key_out;   // calculate.v(9[18:25])
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // calculate.v(3[11:14])
    wire time10ms /* synthesis is_clock=1, SET_AS_NETWORK=time10ms */ ;   // calculate.v(14[9:17])
    
    wire n929, reset_c, key_in_c_3, key_in_c_2, key_in_c_1, key_in_c_0;
    wire [16:0]timecnt;   // calculate.v(13[16:23])
    wire [3:0]scanvalue;   // calculate.v(15[15:24])
    
    wire n8268;
    wire [3:0]flag_Data;   // calculate.v(16[15:24])
    wire [1:0]flag_Cal;   // calculate.v(18[15:23])
    wire [7:0]int_Data0;   // calculate.v(19[15:24])
    
    wire n9152;
    wire [7:0]int_Data1;   // calculate.v(20[15:24])
    
    wire PointTime_c;
    wire [7:0]int_Data;   // calculate.v(22[15:23])
    
    wire key_out_c_3, key_out_c_2, key_out_c_1, key_out_c_0, led_int_Data0_c_3, 
        led_int_Data0_c_2, led_int_Data0_c_1, led_int_Data0_c_0, led_int_Data1_c_3, 
        led_int_Data1_c_2, led_int_Data1_c_1, led_int_Data1_c_0, led_int_Data2_c_3, 
        led_int_Data2_c_0, n32, n4637, n26, n20, n8991, n4, n15, 
        n28, n4549, n9150, time10ms_N_397, n25, n9308, n20_adj_1, 
        n19, n11, n109, n111, n10, n108, n9271, n41, n9148, 
        n35, n9146, n9267, n4_adj_2, n9266, n5861, n10_adj_3, 
        n92, n4491;
    wire [3:0]led_int_Data2_3__N_111;
    
    wire n9140, n9054, n9138, n9136, n15_adj_4, n4608, n8341, 
        n8457, n9134, n3825, n14, n9230, n28_adj_5, n6107, n8978, 
        n4588;
    wire [7:0]int_Data0_7__N_151;
    
    wire n8364, n9128, n8976, n90, n8057, n15_adj_6, n4520, n4567, 
        n9123, n8302, n9268, n96, n5992, n11_adj_7, n6581, n101, 
        n4558, n4609, n3, n9305, n9302, n9296, n1469, n1468, 
        n1467, n1466, n1464, n13, n74, n7, n9122, n89, n103, 
        n78;
    wire [7:0]int_Data1_7__N_351;
    
    wire n22, n15_adj_8, n4490, n4489, n9, n10_adj_9;
    wire [7:0]int_Data0_7__N_183;
    
    wire n29, n11_adj_10, n15_adj_11, n71, n76, n76_adj_12, n97, 
        n9419, n8271, n8263, n1490, n1489, n9418, n9118, n1488, 
        n1487, n1486, n1485, n523, n524, n525, n526, n9030, 
        n9416, n531, n533, n534, n535, n536, n537, n538, n539, 
        n540, n8, n7_adj_13, n6, n4_adj_14, n9113, n3204, n9232, 
        n8259, n8_adj_15, n563, n8395, n8973, n8399, n8400, n8401, 
        n9033, n579, n9380, n9386, n9392, n78_adj_16, n4_adj_17, 
        n8971, n94, led_int_Data2_3__N_109, n8354;
    wire [3:0]led_int_Data2_3__N_67;
    
    wire n9108, n5, n145, n8305, n91, led_int_Data1_3__N_385, n9398, 
        n731, n9404, n9410, n4148, n4564, n744, n8349, n757, 
        n8968, n4645, n34, n770, n783, n1524, n796, n10_adj_18, 
        n9116, n4607, n22_adj_19, n9018, n9106, n9415, n6101, 
        n6099, n8262, n14_adj_20, n8_adj_21, n8386, n8254, n8253, 
        n854, n4459, n9414, n858, n9412, n862, n864, n9338, 
        n9341, n9344, n5850, n874, n17, n9_adj_22;
    wire [3:0]led_int_Data1_3__N_381;
    wire [3:0]led_int_Data0_3__N_388;
    wire [3:0]led_int_Data1_3__N_63;
    wire [3:0]led_int_Data0_3__N_59;
    
    wire n1512, n1511, n9102, n9048, n9411, n9409, n4638, n9408, 
        n9406, n9405, n9403, n8680, n6_adj_23, n3205, n4586, n3206, 
        n1207, n6_adj_24, n1208, n9016, n9068, n19_adj_25, n6093, 
        n5887, n104, n9_adj_26, n1491, n1480, n70, n31, n9241, 
        n1298, n1299, n1300, n1305, n1311, n1317, n1323, n1329, 
        n1556, n102, n82, n9_adj_27, n124, n5883, n100, n97_adj_28, 
        n16, n9280, n29_adj_29, n8313, n32_adj_30, n4546, n9277, 
        n91_adj_31, n104_adj_32, n4492, n4543, n8315, n78_adj_33, 
        n9402, n4561, n9021, n5880, n9400, n9399, n9397, n9396, 
        n85, n79, n1701, n9374, n9326, n29_adj_34, n9082, n8177, 
        n9239, n17_adj_35, n75, n21, n8336, n9100, n9092, n4_adj_36, 
        n8064, n8241, n19_adj_37, n4572, n9098, n4783, n38, n8_adj_38, 
        n9265, n9394, n5957, n6225, n5835, n9256, n16_adj_39, 
        n9259, n4292, n5955, n5874, n9393, n9391, n3504, n8982, 
        n8964, n15_adj_40, n3830, n3842, n13_adj_41, n9012, n22_adj_42, 
        n169, n73, n112, n9274, n5953, n92_adj_43, n15_adj_44, 
        n8173, n15_adj_45, n9008, n9390, n11_adj_46, n9_adj_47, 
        n9285, n9388, n9290, n4149, n9387, n8999, n2, n4_adj_48, 
        n97_adj_49, n12, n9317, n31_adj_50, n6214, n82_adj_51, n8360, 
        n8250, n66, n9385, n72, n74_adj_52, n115, n67, n68, 
        n9262, n93, n15_adj_53, n79_adj_54, n55, n8348, n9004, 
        n47, n9104, n9022, n12_adj_55, n9_adj_56, n69, n70_adj_57, 
        n9234, n43, n10_adj_58, n67_adj_59, n82_adj_60, n52, n8498, 
        n88, n4_adj_61, n8176, n9384, n9382, n8_adj_62, n9381, 
        n9028, n75_adj_63, n8078, n9379, n64, n9238, n4_adj_64, 
        n4_adj_65, n66_adj_66, n6_adj_67, n4_adj_68, n21_adj_69, n4_adj_70, 
        n87, n12_adj_71, n9378, n8318, n94_adj_72, n15_adj_73, n14_adj_74, 
        n9376, n106, n4651, n22_adj_75, n4_adj_76, n9375, n9373, 
        n8_adj_77, n67_adj_78, n8393, n9035, n9112, n10_adj_79, 
        n9284, n106_adj_80, n15_adj_81, n9031, n9_adj_82, n8168, 
        n6052, n14_adj_83, n9372, n3_adj_84, n4_adj_85, n9370, n6_adj_86, 
        n9369, n9311, n4535, n9368, n7960, n95, n15_adj_87, n4_adj_88, 
        n6191, n7_adj_89, n8326, n8712, n6189, n6167, n4_adj_90, 
        n16_adj_91, n66_adj_92, n5_adj_93, n4_adj_94, n6_adj_95, n4644, 
        n4_adj_96, n4_adj_97, n6042, n6_adj_98, n9413, n8504, n6038, 
        n4587, n6_adj_99, n4_adj_100, n10_adj_101, n5869, n15_adj_102, 
        n9229, n5812, n4293, n9365, n99, n9362, n9359, n9282, 
        n4712, n8340, n8317, n8444, n9299, n8986, n68_adj_103, 
        n72_adj_104, n73_adj_105, n8506, n15_adj_106, n14_adj_107, 
        n8979, n4698, n9320, n4554, n9248, n7946, n9366, n8164, 
        n15_adj_108, n9356, n9353, n148, n6181, n4245, n87_adj_109, 
        n8963, n9251, n8961, n5_adj_110, n9350, n4789, n9281, 
        n8993, n9347, n79_adj_111, n22_adj_112, n8959, n9364, n15_adj_113, 
        n14_adj_114, n6026, n5926, n6089, n3435, n4686, n9013, 
        n11_adj_115, n4684, n5829, n4495, n4682, n5921, n14_adj_116, 
        n4639, n6_adj_117, n9407, n4681, n8167, n4680, n4679, 
        n5843, n6314, n3967, n9363, n3759, n3722, n5859, n6171, 
        n4244, n5856, n90_adj_118, n15_adj_119, n3758, n13_adj_120, 
        n9243, n10_adj_121, n18, n5854, n8310, n9401, n8229, n6020, 
        n77, n28_adj_122, n69_adj_123, n4_adj_124, n8071, n21_adj_125, 
        n9361, n9236, n40, n8159, n5916, n9007, n9283, n8_adj_126, 
        n3513, n49, n4787, n9360, n79_adj_127, n3724, n7953, n9005, 
        n100_adj_128, n4_adj_129, n8950, n9358, n22_adj_130, n84, 
        n9357, n80, n9355, n83, n84_adj_131, n8335, n21_adj_132, 
        n15_adj_133, n55_adj_134, n9354, n4_adj_135, n7_adj_136, n5797, 
        n6_adj_137, n12_adj_138, n8988, n4_adj_139, n7942, n4391, 
        n6150, n24, n9_adj_140, n3187, n9253, n4_adj_141, n38_adj_142, 
        n5826, n85_adj_143, n9383, n34_adj_144, n9286, n68_adj_145, 
        n4548, n9389, n22_adj_146, n9377, n8225, n92_adj_147, n50, 
        n86, n9002, n19_adj_148, n9352, n9395, n4_adj_149, n9351, 
        n4555, n49_adj_150, n5913, n28_adj_151, n8339, n4_adj_152, 
        n9349, n9348, n4540, n4355, n9346, n9345, n3757, n5841, 
        n3721, n9343, n127, n4090, n9342, n8158, n9323, n9340, 
        n9339, n5999, n9337, n9051, n9336, n18_adj_153, n6141, 
        n3725, n9335, n1, n41_adj_154, n8480, n8477, n11_adj_155, 
        n1_adj_156, n4067, n4066, n8345, n5839, n6133, n6368, 
        n3760, n8473, n8343, n9010, n8468, n6123, n8467, n3723, 
        n5820, n8464, n8228, n8458, n5795, n9242, n8220, n5837, 
        n9333, n8452, n9019, n4_adj_157, n9245, n9006, n9003, 
        n9332, n9065, n9064, n4_adj_158, n8441, n8598, n8439, 
        n121, n4475, n58, n4473, n4471, n25_adj_159, n8980, n8398, 
        n8352, n8388, n9330, n6111, n9060, n4464, n9124, n9_adj_160, 
        n4462, n9246, n9329, n4_adj_161, n8146, n8437, n8216, 
        n8005, n4_adj_162, n4_adj_163, n6_adj_164, n7911, n6_adj_165, 
        n8001, n8435, n8219, n4_adj_166, n8_adj_167, n7920, n8050, 
        n8211, n7938, n8433, n8155, n9063, n8004, n8207, n4_adj_168, 
        n14_adj_169, n10_adj_170, n7941, n7933, n8429, n8290, n8427, 
        n8210, n7996, n8202, n6_adj_171, n8425, n8201, n8955, 
        n8286, n7992, n7929, n8189, n8134, n8127, n8_adj_172, 
        n8120, n7995, n8_adj_173, n7987, n8289, n8953, n8113, 
        n8106, n7983, n9250, n8198, n8099, n10_adj_174, n8_adj_175, 
        n7986, n8281, n8092, n7932, n8948, n9080, n8277, n7924, 
        n8085, n8300, n7923, n4_adj_176, n9327, n4_adj_177, n4_adj_178, 
        n9325, n9045, n1_adj_179, n8642, n9324, n9072, n10_adj_180, 
        n8_adj_181, pwr, n9371, n8280, n8272, n8590, n6_adj_182, 
        n4_adj_183, n4_adj_184, n9287, n1_adj_185, n3_adj_186, n6_adj_187, 
        n9321, n9417, n9319, n9142, n19_adj_188, n24_adj_189, n25_adj_190, 
        n8744, n9318, n9316, n9315, n9314, n9312, n9040, n9310, 
        n9309, n9307, n9306, n9304, n9303, n9301, n4_adj_191, 
        n9300, n9017, n9298, n9297, n9295, n9294, n9293, n9291, 
        n9289, n9288, n9057, n9279, n9263, n9027, n9278, n9260, 
        n9276, n1_adj_192, n9257, n9275, n16_adj_193, n15_adj_194, 
        n9254, n8996, n9219, n4_adj_195, n9218, n9273, n9205, 
        n9203, n9202, n9200, n9198, n9015, n1_adj_196, n4_adj_197, 
        n9272, n9086, n9192, n9188, n9227, n9233, n9180, n9178, 
        n9217, n9172, n9211, n9168, n4_adj_198, n12_adj_199, n9164, 
        n9162, n9269, n9154;
    
    AND2 mult_119_i86 (.O(n127), .I0(int_Data1[2]), .I1(int_Data0[5]));
    AND2 i6695 (.O(n9345), .I0(n1300), .I1(n1485));
    AND2 mult_119_i98 (.O(n145), .I0(int_Data1[0]), .I1(int_Data0[6]));
    AND5 i4 (.O(n9003), .I0(n5850), .I1(n5820), .I2(n15_adj_4), .I3(n9002), 
         .I4(n15_adj_113));
    AND2 mult_119_i100 (.O(n148), .I0(int_Data1[1]), .I1(int_Data0[6]));
    OR2 i5624 (.O(n8262), .I0(n4_adj_76), .I1(n73));
    AND2 mult_119_i114 (.O(n169), .I0(int_Data1[0]), .I1(int_Data0[7]));
    OR2 i977 (.O(n6_adj_117), .I0(int_Data[2]), .I1(int_Data[1]));
    XOR2 i5604 (.O(n579), .I0(n25_adj_159), .I1(n5));
    OR2 i5625 (.O(n6_adj_67), .I0(n8259), .I1(n8263));
    DFFCR int_Data1_i0_i2 (.Q(int_Data1[2]), .D(n4645), .CLK(time10ms), 
          .CE(n4679), .R(reset_c));   // calculate.v(55[13] 193[16])
    DFFCR flag_Data_i0 (.Q(flag_Data[0]), .D(n8590), .CLK(time10ms), .CE(n4682), 
          .R(reset_c));   // calculate.v(55[13] 193[16])
    XOR2 i5557 (.O(n3725), .I0(n28_adj_5), .I1(n8_adj_38));
    OR2 i6483 (.O(n9128), .I0(n9005), .I1(n9068));
    DFFCR int_Data1_i0_i1 (.Q(int_Data1[1]), .D(n4639), .CLK(time10ms), 
          .CE(n4679), .R(reset_c));   // calculate.v(55[13] 193[16])
    DFFC key_out_i0_i1 (.Q(key_out_c_0), .D(scanvalue[0]), .CLK(time10ms), 
         .CE(reset_c));   // calculate.v(55[13] 193[16])
    DFFCR led_int_Data2_i1 (.Q(led_int_Data2_c_0), .D(led_int_Data2_3__N_67[0]), 
          .CLK(time10ms), .CE(n4686), .R(reset_c));   // calculate.v(55[13] 193[16])
    DFFCS PointTime_223 (.Q(PointTime_c), .D(n8364), .CLK(time10ms), .CE(n19_adj_188), 
          .S(reset_c));   // calculate.v(55[13] 193[16])
    DFFCR int_Data0_i0_i0 (.Q(int_Data0[0]), .D(n8712), .CLK(time10ms), 
          .CE(n4679), .R(reset_c));   // calculate.v(55[13] 193[16])
    DFFR led_int_Data1_i1 (.Q(led_int_Data1_c_0), .D(led_int_Data1_3__N_63[0]), 
         .CLK(clk_c), .R(reset_c));   // calculate.v(204[13] 242[16])
    DFFR led_int_Data0_i1 (.Q(led_int_Data0_c_0), .D(led_int_Data0_3__N_388[0]), 
         .CLK(clk_c), .R(reset_c));   // calculate.v(204[13] 242[16])
    OR2 i1126 (.O(n4_adj_88), .I0(n3513), .I1(n4149));
    AND2 i2199 (.O(n4783), .I0(n11_adj_46), .I1(n11_adj_115));
    XOR2 i5518 (.O(n3760), .I0(n31_adj_50), .I1(n11_adj_155));
    XOR2 i1035 (.O(n858), .I0(int_Data[1]), .I1(n4355));
    XOR2 i1_adj_1 (.O(n4475), .I0(n6171), .I1(n8437));
    OR2 i6696 (.O(n9346), .I0(n9345), .I1(n9344));
    OR2 i1_adj_2 (.O(n79), .I0(n1208), .I1(flag_Data[0]));
    DFFR scanvalue_FSM_i0 (.Q(scanvalue[3]), .D(scanvalue[2]), .CLK(time10ms), 
         .R(reset_c));   // calculate.v(57[17] 63[24])
    DFFR timecnt_941_942__i15 (.Q(timecnt[14]), .D(n83), .CLK(clk_c), 
         .R(reset_c)) /* synthesis syn_use_carry_chain=1 */ ;   // calculate.v(36[23:32])
    AND2 i5626 (.O(n8263), .I0(n8262), .I1(n3724));
    DFFR timecnt_941_942__i14 (.Q(timecnt[13]), .D(n84_adj_131), .CLK(clk_c), 
         .R(reset_c)) /* synthesis syn_use_carry_chain=1 */ ;   // calculate.v(36[23:32])
    DFFR timecnt_941_942__i13 (.Q(timecnt[12]), .D(n85_adj_143), .CLK(clk_c), 
         .R(reset_c)) /* synthesis syn_use_carry_chain=1 */ ;   // calculate.v(36[23:32])
    DFFR timecnt_941_942__i12 (.Q(timecnt[11]), .D(n86), .CLK(clk_c), 
         .R(reset_c)) /* synthesis syn_use_carry_chain=1 */ ;   // calculate.v(36[23:32])
    DFFR timecnt_941_942__i11 (.Q(timecnt[10]), .D(n87), .CLK(clk_c), 
         .R(reset_c)) /* synthesis syn_use_carry_chain=1 */ ;   // calculate.v(36[23:32])
    DFFR timecnt_941_942__i10 (.Q(timecnt[9]), .D(n88), .CLK(clk_c), .R(reset_c)) /* synthesis syn_use_carry_chain=1 */ ;   // calculate.v(36[23:32])
    DFFR timecnt_941_942__i9 (.Q(timecnt[8]), .D(n89), .CLK(clk_c), .R(reset_c)) /* synthesis syn_use_carry_chain=1 */ ;   // calculate.v(36[23:32])
    DFFR timecnt_941_942__i8 (.Q(timecnt[7]), .D(n90), .CLK(clk_c), .R(reset_c)) /* synthesis syn_use_carry_chain=1 */ ;   // calculate.v(36[23:32])
    INV i1256 (.O(n3842), .I0(flag_Data[1]));
    DFFR timecnt_941_942__i1 (.Q(timecnt[0]), .D(n80), .CLK(clk_c), .R(reset_c)) /* synthesis syn_use_carry_chain=1 */ ;   // calculate.v(36[23:32])
    AND2 i1_adj_3 (.O(n4608), .I0(n70_adj_57), .I1(n4607));
    DFFR timecnt_941_942__i7 (.Q(timecnt[6]), .D(n91), .CLK(clk_c), .R(reset_c)) /* synthesis syn_use_carry_chain=1 */ ;   // calculate.v(36[23:32])
    DFFR timecnt_941_942__i6 (.Q(timecnt[5]), .D(n92_adj_43), .CLK(clk_c), 
         .R(reset_c)) /* synthesis syn_use_carry_chain=1 */ ;   // calculate.v(36[23:32])
    OR2 i3694 (.O(n6314), .I0(n6171), .I1(n535));
    AND2 i5319 (.O(n7942), .I0(n7941), .I1(int_Data0[3]));
    DFFCR int_Data1_i0_i0 (.Q(int_Data1[0]), .D(n4609), .CLK(time10ms), 
          .CE(n4679), .R(reset_c));   // calculate.v(55[13] 193[16])
    DFFR timecnt_941_942__i5 (.Q(timecnt[4]), .D(n93), .CLK(clk_c), .R(reset_c)) /* synthesis syn_use_carry_chain=1 */ ;   // calculate.v(36[23:32])
    AND2 i6698 (.O(n9348), .I0(n1300), .I1(n1486));
    DFFR timecnt_941_942__i4 (.Q(timecnt[3]), .D(n94_adj_72), .CLK(clk_c), 
         .R(reset_c)) /* synthesis syn_use_carry_chain=1 */ ;   // calculate.v(36[23:32])
    DFFR timecnt_941_942__i3 (.Q(timecnt[2]), .D(n95), .CLK(clk_c), .R(reset_c)) /* synthesis syn_use_carry_chain=1 */ ;   // calculate.v(36[23:32])
    DFFR timecnt_941_942__i2 (.Q(timecnt[1]), .D(n96), .CLK(clk_c), .R(reset_c)) /* synthesis syn_use_carry_chain=1 */ ;   // calculate.v(36[23:32])
    DFFCR flag_Cal_i0_i0 (.Q(flag_Cal[0]), .D(n5856), .CLK(time10ms), 
          .CE(n1480), .R(reset_c));   // calculate.v(55[13] 193[16])
    OR2 i6759 (.O(n9409), .I0(n9408), .I1(n9407));
    AND3 i2 (.O(n8313), .I0(n9057), .I1(int_Data1[0]), .I2(n5887));
    XOR2 i5321 (.O(n526), .I0(n8_adj_173), .I1(int_Data0[4]));
    INV i30 (.O(n4586), .I0(n97));
    XOR2 i2_adj_4 (.O(n8395), .I0(n4_adj_90), .I1(n145));
    OR2 i1_adj_5 (.O(n4651), .I0(n8300), .I1(n8961));
    OR2 key_in_3__I_0_239_i10 (.O(n10_adj_121), .I0(key_out_c_3), .I1(key_out_c_2));
    OR2 i6485 (.O(n9068), .I0(n9122), .I1(n19_adj_25));
    AND2 i1_adj_6 (.O(n97), .I0(n6167), .I1(n15_adj_113));
    AND2 i6721 (.O(n9371), .I0(n4491), .I1(n9346));
    AND3 i2_adj_7 (.O(n8310), .I0(n50), .I1(n92_adj_147), .I2(n4_adj_94));
    OR2 i1_adj_8 (.O(int_Data1_7__N_351[3]), .I0(n66), .I1(n92));
    AND2 i1_adj_9 (.O(n8590), .I0(n9370), .I1(n5795));
    OR2 i6699 (.O(n9349), .I0(n9348), .I1(n9347));
    AND2 i5371 (.O(n7996), .I0(n7995), .I1(int_Data0[2]));
    AND2 i6701 (.O(n9351), .I0(n1300), .I1(n1487));
    AND2 i1_adj_10 (.O(n4638), .I0(n75), .I1(n4637));
    XOR2 i1_adj_11 (.O(n4462), .I0(n6099), .I1(n8441));
    AND2 i3297 (.O(n1468), .I0(n5869), .I1(n9388));
    AND3 i6718 (.O(n9368), .I0(n5921), .I1(n3842), .I2(n1701));
    OR2 i1_adj_12 (.O(n15_adj_73), .I0(n14_adj_74), .I1(n11_adj_115));
    OR2 i3216 (.O(n5797), .I0(n783), .I1(n770));
    AND2 i1_adj_13 (.O(n8999), .I0(n38_adj_142), .I1(n10));
    OR2 equal_433_i17 (.O(n17), .I0(n16_adj_39), .I1(n14_adj_20));
    OR2 i1_adj_14 (.O(n75), .I0(n69), .I1(n92));
    AND2 i1_adj_15 (.O(n94), .I0(n15_adj_102), .I1(n15_adj_108));
    OR2 i6702 (.O(n9352), .I0(n9351), .I1(n9350));
    AND2 i3300 (.O(n1469), .I0(n5869), .I1(n9394));
    AND2 i6704 (.O(n9354), .I0(n1300), .I1(n1488));
    OR2 i1_adj_16 (.O(n74_adj_52), .I0(n1701), .I1(n1208));
    OR2 key_in_3__I_0_241_i15 (.O(n15_adj_119), .I0(n14), .I1(n11_adj_10));
    OR2 i6705 (.O(n9355), .I0(n9354), .I1(n9353));
    AND2 i1_adj_17 (.O(n3), .I0(n15_adj_11), .I1(n15_adj_113));
    AND2 i3339 (.O(n5921), .I0(n9232), .I1(n15_adj_53));
    OR2 i3571 (.O(n6171), .I0(n6099), .I1(n536));
    OR2 key_in_3__I_0_238_i15 (.O(n15_adj_4), .I0(n14), .I1(n11_adj_7));
    INV i554 (.O(n1511), .I0(led_int_Data1_3__N_385));
    OR2 i1_adj_18 (.O(n72), .I0(n68), .I1(n92));
    OR2 i1_adj_19 (.O(n9112), .I0(n4_adj_2), .I1(n8964));
    AND2 i5631 (.O(n8268), .I0(n6_adj_67), .I1(n97_adj_49));
    AND2 i1_adj_20 (.O(n4644), .I0(n72), .I1(n4586));
    INV i6429 (.O(n9019), .I0(n9068));
    OR2 i5632 (.O(n8271), .I0(n6_adj_67), .I1(n97_adj_49));
    AND4 i3 (.O(n9004), .I0(n9002), .I1(n5992), .I2(n3), .I3(n5926));
    OR2 key_in_3__I_0_239_i15 (.O(n15_adj_6), .I0(n14_adj_114), .I1(n11_adj_10));
    INV i1135 (.O(n10), .I0(key_in_c_1));
    OR2 i1_adj_21 (.O(n9015), .I0(n9013), .I1(key_in_c_2));
    INV i292 (.O(n563), .I0(n531));
    XOR2 i1_adj_22 (.O(n4464), .I0(n5861), .I1(n8429));
    OR2 i1_adj_23 (.O(n9017), .I0(n9016), .I1(n9_adj_22));
    AND2 i6707 (.O(n9357), .I0(n1300), .I1(n1489));
    OR2 i3630 (.O(n6167), .I0(n6189), .I1(n11_adj_10));
    XOR2 i6 (.O(n8393), .I0(n12_adj_199), .I1(n11));
    AND2 i5431 (.O(n8057), .I0(n8050), .I1(timecnt[2]));
    OR2 i6708 (.O(n9358), .I0(n9357), .I1(n9356));
    OR2 i1_adj_24 (.O(n4_adj_48), .I0(n16), .I1(n22_adj_42));
    AND2 i6710 (.O(n9360), .I0(n1300), .I1(n1490));
    OR2 i6711 (.O(n9361), .I0(n9360), .I1(n9359));
    OR2 key_in_3__I_0_237_i11 (.O(n11_adj_7), .I0(n10_adj_121), .I1(n16_adj_39));
    AND2 i6713 (.O(n9363), .I0(n1300), .I1(n1491));
    OR2 i1_adj_25 (.O(n21_adj_132), .I0(n9_adj_140), .I1(key_in_c_2));
    AND2 i1_adj_26 (.O(n55), .I0(n9021), .I1(n6_adj_24));
    AND2 i3271 (.O(n5859), .I0(n14_adj_114), .I1(n14));
    AND3 i1_adj_27 (.O(n8973), .I0(n8955), .I1(n5837), .I2(n5835));
    INV i1027 (.O(n7_adj_136), .I0(int_Data[3]));
    AND2 i6469 (.O(n9113), .I0(n9112), .I1(n8458));
    OR2 i6714 (.O(n9364), .I0(n9363), .I1(n9362));
    AND2 i6633 (.O(n9283), .I0(n9256), .I1(n5921));
    OR2 key_in_3__I_0_238_i14 (.O(n14), .I0(n13_adj_120), .I1(n9013));
    AND2 i6716 (.O(n9366), .I0(flag_Data[1]), .I1(int_Data0[2]));
    OR2 i6717 (.O(int_Data0_7__N_151[2]), .I0(n9366), .I1(n9365));
    OR2 key_in_3__I_0_240_i9 (.O(n16), .I0(n19), .I1(key_out_c_0));
    XOR2 i5421 (.O(n79_adj_127), .I0(timecnt[0]), .I1(timecnt[1]));
    OR2 key_in_3__I_0_239_i11 (.O(n11_adj_10), .I0(n10_adj_121), .I1(n16));
    AND2 i5576 (.O(n8207), .I0(n4_adj_183), .I1(n76));
    OR2 i5633 (.O(n8_adj_62), .I0(n8268), .I1(n8272));
    OR2 i5577 (.O(n8210), .I0(n4_adj_183), .I1(n76));
    AND2 i6719 (.O(n9369), .I0(flag_Data[1]), .I1(n9285));
    OR2 i6720 (.O(n9370), .I0(n9369), .I1(n9368));
    OR2 i3577 (.O(n5913), .I0(n6225), .I1(n14));
    DFFS scanvalue_FSM_i3 (.Q(scanvalue[0]), .D(scanvalue[3]), .CLK(time10ms), 
         .S(reset_c));   // calculate.v(57[17] 63[24])
    OR2 i6626 (.O(n9276), .I0(n9275), .I1(n9274));
    OR2 i5578 (.O(n6_adj_182), .I0(n8207), .I1(n8211));
    OR2 key_in_3__I_0_240_i15 (.O(n15_adj_133), .I0(n14_adj_107), .I1(n11_adj_10));
    AND2 i6761 (.O(n9411), .I0(n1298), .I1(n9035));
    AND2 i1_adj_28 (.O(n67_adj_78), .I0(n66_adj_66), .I1(n9_adj_82));
    AND2 i3408 (.O(n5992), .I0(n15_adj_133), .I1(n15_adj_4));
    OR2 key_in_3__I_0_237_i9 (.O(n16_adj_39), .I0(key_out_c_1), .I1(n20_adj_1));
    OR2 equal_936_i14 (.O(n7_adj_89), .I0(flag_Data[1]), .I1(led_int_Data2_3__N_111[1]));
    OR2 i3407 (.O(n9104), .I0(n8968), .I1(n4_adj_184));
    AND2 i5579 (.O(n8211), .I0(n8210), .I1(n3759));
    AND2 i1_adj_29 (.O(n4_adj_2), .I0(n9048), .I1(n12_adj_71));
    AND2 i5634 (.O(n8272), .I0(n8271), .I1(n3723));
    AND2 i6647 (.O(n9297), .I0(key_out_c_2), .I1(n115));
    OR3 i3578 (.O(n5916), .I0(n9086), .I1(n13), .I2(n11_adj_10));
    XOR2 i5442 (.O(n76_adj_12), .I0(n8064), .I1(timecnt[4]));
    OR2 key_in_3__I_0_236_i15 (.O(n15_adj_8), .I0(n14_adj_114), .I1(n11_adj_7));
    AND2 i1_adj_30 (.O(n32), .I0(n9015), .I1(key_in_c_3));
    AND2 i6722 (.O(n9372), .I0(n1299), .I1(n533));
    OR2 equal_936_i22 (.O(n22), .I0(n21), .I1(n19_adj_25));
    XOR2 i5449 (.O(n75_adj_63), .I0(n8071), .I1(timecnt[5]));
    AND2 i3579 (.O(n6181), .I0(n9008), .I1(n15_adj_73));
    OR2 equal_412_i20 (.O(n13_adj_120), .I0(key_in_c_3), .I1(n9_adj_27));
    AND2 i3269 (.O(n5850), .I0(n15_adj_6), .I1(n15_adj_11));
    AND2 i6462 (.O(n3205), .I0(n9104), .I1(n8468));
    XOR2 i1_adj_31 (.O(n8437), .I0(n10_adj_170), .I1(int_Data0[5]));
    OR2 equal_425_i21 (.O(n21), .I0(n13), .I1(n10));
    AND2 i1_adj_32 (.O(n64), .I0(n8953), .I1(n47));
    AND2 i1_adj_33 (.O(n15), .I0(key_in_c_0), .I1(key_in_c_1));
    AND2 i1_adj_34 (.O(n26), .I0(key_out_c_0), .I1(key_out_c_1));
    OR2 equal_412_i21 (.O(n21_adj_125), .I0(n13_adj_120), .I1(key_in_c_1));
    OR2 i6723 (.O(n9373), .I0(n9372), .I1(n9371));
    AND4 i6628 (.O(n9278), .I0(n4543), .I1(key_out_c_3), .I2(key_in_c_3), 
         .I3(n8986));
    AND2 i6630 (.O(n9280), .I0(led_int_Data2_3__N_109), .I1(n9072));
    OR2 i1_adj_35 (.O(n66_adj_66), .I0(n79_adj_54), .I1(n55));
    INV i849 (.O(n1524), .I0(n731));
    AND2 i6725 (.O(n9375), .I0(n1298), .I1(n523));
    AND4 i6627 (.O(n9277), .I0(flag_Data[0]), .I1(n4540), .I2(n29_adj_29), 
         .I3(n32_adj_30));
    OR2 equal_424_i22 (.O(n22_adj_19), .I0(n21), .I1(n19_adj_148));
    OR2 i6488 (.O(n9134), .I0(n5859), .I1(n11_adj_10));
    OR2 i3279 (.O(n5861), .I0(n540), .I1(n539));
    OR2 equal_412_i22 (.O(n22_adj_112), .I0(n21_adj_125), .I1(n19_adj_25));
    AND3 i6490 (.O(n9136), .I0(n8991), .I1(n15_adj_4), .I2(n15_adj_108));
    AND2 i1_adj_36 (.O(n6_adj_98), .I0(flag_Data[0]), .I1(n29_adj_29));
    INV i24 (.O(n4637), .I0(n78_adj_16));
    AND2 i1_adj_37 (.O(n104_adj_32), .I0(n9276), .I1(n10));
    AND2 i5337 (.O(n7960), .I0(n7953), .I1(int_Data0[6]));
    OR2 i6726 (.O(n9376), .I0(n9375), .I1(n9374));
    AND2 i6728 (.O(n9378), .I0(n1299), .I1(n534));
    OR2 i6729 (.O(n9379), .I0(n9378), .I1(n9377));
    AND2 i3218 (.O(n83), .I0(n29), .I1(n66_adj_92));
    AND2 i3430 (.O(n6225), .I0(n11_adj_7), .I1(n11_adj_115));
    AND2 i6715 (.O(n9365), .I0(n3842), .I1(led_int_Data2_3__N_111[1]));
    AND2 i6712 (.O(n9362), .I0(n4490), .I1(n579));
    INV i3231 (.O(n5812), .I0(n757));
    AND2 i6709 (.O(n9359), .I0(n4490), .I1(n8401));
    OR2 equal_421_i22 (.O(n22_adj_146), .I0(n21_adj_125), .I1(n19_adj_148));
    DFFR scanvalue_FSM_i2 (.Q(scanvalue[1]), .D(scanvalue[0]), .CLK(time10ms), 
         .R(reset_c));   // calculate.v(57[17] 63[24])
    DFFR scanvalue_FSM_i1 (.Q(scanvalue[2]), .D(scanvalue[1]), .CLK(time10ms), 
         .R(reset_c));   // calculate.v(57[17] 63[24])
    DFFCR int_Data__i8 (.Q(int_Data[7]), .D(n1466), .CLK(time10ms), .CE(n4698), 
          .R(reset_c));   // calculate.v(55[13] 193[16])
    DFFCR int_Data__i7 (.Q(int_Data[6]), .D(n1467), .CLK(time10ms), .CE(n4698), 
          .R(reset_c));   // calculate.v(55[13] 193[16])
    DFFR led_int_Data0_i4 (.Q(led_int_Data0_c_3), .D(led_int_Data0_3__N_59[3]), 
         .CLK(clk_c), .R(reset_c));   // calculate.v(204[13] 242[16])
    DFFR led_int_Data0_i3 (.Q(led_int_Data0_c_2), .D(led_int_Data0_3__N_59[2]), 
         .CLK(clk_c), .R(reset_c));   // calculate.v(204[13] 242[16])
    DFFCR int_Data__i6 (.Q(int_Data[5]), .D(n1468), .CLK(time10ms), .CE(n4698), 
          .R(reset_c));   // calculate.v(55[13] 193[16])
    DFFCR int_Data__i5 (.Q(int_Data[4]), .D(n1469), .CLK(time10ms), .CE(n4698), 
          .R(reset_c));   // calculate.v(55[13] 193[16])
    DFFCR int_Data__i4 (.Q(int_Data[3]), .D(n9295), .CLK(time10ms), .CE(n4698), 
          .R(reset_c));   // calculate.v(55[13] 193[16])
    DFFR led_int_Data0_i2 (.Q(led_int_Data0_c_1), .D(led_int_Data0_3__N_59[1]), 
         .CLK(clk_c), .R(reset_c));   // calculate.v(204[13] 242[16])
    DFFCR int_Data__i3 (.Q(int_Data[2]), .D(n9301), .CLK(time10ms), .CE(n4698), 
          .R(reset_c));   // calculate.v(55[13] 193[16])
    DFFCR int_Data__i2 (.Q(int_Data[1]), .D(n9304), .CLK(time10ms), .CE(n4698), 
          .R(reset_c));   // calculate.v(55[13] 193[16])
    DFFCR flag_Cal_i0_i1 (.Q(flag_Cal[1]), .D(n5826), .CLK(time10ms), 
          .CE(n1480), .R(reset_c));   // calculate.v(55[13] 193[16])
    OR2 i6629 (.O(n9279), .I0(n9278), .I1(n9277));
    OR2 equal_421_i19 (.O(n19_adj_148), .I0(n18), .I1(key_out_c_2));
    OR5 i4_adj_38 (.O(n4489), .I0(key_out_c_2), .I1(flag_Cal[0]), .I2(n4558), 
        .I3(n9_adj_47), .I4(n1));
    OR2 i1_adj_39 (.O(n100), .I0(n91_adj_31), .I1(n8315));
    OR2 i3436 (.O(n5837), .I0(n6026), .I1(n22_adj_146));
    AND2 i3344 (.O(n5926), .I0(n15_adj_6), .I1(n15_adj_106));
    OR2 i1_adj_40 (.O(n97_adj_28), .I0(n84), .I1(n82));
    AND2 i6706 (.O(n9356), .I0(n4490), .I1(n8400));
    AND2 i1_adj_41 (.O(n91_adj_31), .I0(n9298), .I1(n19));
    AND2 i5323 (.O(n7946), .I0(n8_adj_173), .I1(int_Data0[4]));
    AND2 i6703 (.O(n9353), .I0(n4490), .I1(n8399));
    AND2 i6700 (.O(n9350), .I0(n4490), .I1(n8398));
    AND2 i6697 (.O(n9347), .I0(n4490), .I1(n8395));
    OR2 i3587 (.O(n5953), .I0(n6189), .I1(n11_adj_7));
    OR2 i1_adj_42 (.O(n9018), .I0(n9016), .I1(n8973));
    OR2 i1_adj_43 (.O(n9006), .I0(n9005), .I1(n22_adj_112));
    AND2 i3346 (.O(n6141), .I0(n14_adj_107), .I1(n14));
    OR2 equal_413_i14 (.O(n14_adj_83), .I0(flag_Data[1]), .I1(flag_Data[0]));
    INV i6579 (.O(n9229), .I0(n4572));
    OR2 equal_934_i18 (.O(n18_adj_153), .I0(n31), .I1(key_out_c_3));
    OR2 i1_adj_44 (.O(n15_adj_113), .I0(n14_adj_114), .I1(n11_adj_115));
    AND2 i1_adj_45 (.O(n78_adj_16), .I0(n3), .I1(n6214));
    INV i5824 (.O(n8464), .I0(n12_adj_71));
    OR2 i1_adj_46 (.O(n9005), .I0(n9_adj_47), .I1(flag_Data[0]));
    AND2 i2_adj_47 (.O(n4391), .I0(n4_adj_68), .I1(n6_adj_86));
    OR2 i2201 (.O(n5795), .I0(n4783), .I1(n14_adj_74));
    XOR2 i2_adj_48 (.O(led_int_Data0_3__N_388[3]), .I0(n4_adj_139), .I1(n4_adj_88));
    OR2 i6762 (.O(n9412), .I0(n9411), .I1(n9410));
    XOR2 i5456 (.O(n74), .I0(n8078), .I1(timecnt[6]));
    AND2 i5639 (.O(n8277), .I0(n8_adj_62), .I1(n121));
    OR2 equal_418_i21 (.O(n21_adj_69), .I0(n13), .I1(key_in_c_1));
    OR2 i1_adj_49 (.O(n4_adj_124), .I0(n4520), .I1(n796));
    OR2 i6440 (.O(n8982), .I0(n9080), .I1(n14_adj_114));
    AND2 i6731 (.O(n9381), .I0(n1298), .I1(n524));
    AND3 i6492 (.O(n9138), .I0(n15_adj_102), .I1(n9134), .I2(n6150));
    OR2 i5640 (.O(n8280), .I0(n8_adj_62), .I1(n121));
    AND2 i1_adj_50 (.O(n4682), .I0(n4680), .I1(n4681));
    XOR2 i5435 (.O(n77), .I0(n8057), .I1(timecnt[3]));
    OR2 i5641 (.O(n10_adj_58), .I0(n8277), .I1(n8281));
    AND5 i3_adj_51 (.O(n16_adj_193), .I0(n4_adj_96), .I1(n15_adj_194), 
         .I2(n8477), .I3(int_Data[6]), .I4(n5957));
    AND2 i6694 (.O(n9344), .I0(n4490), .I1(n8393));
    OR2 key_in_3__I_0_243_i15 (.O(n15_adj_106), .I0(n14_adj_107), .I1(n11_adj_115));
    AND2 i6456 (.O(n9098), .I0(n5829), .I1(n6107));
    AND2 i6691 (.O(n9341), .I0(n5812), .I1(n858));
    DFFC time10ms_215 (.Q(time10ms), .D(time10ms_N_397), .CLK(clk_c), 
         .CE(reset_c));   // calculate.v(31[14] 36[33])
    AND2 i6450 (.O(n9092), .I0(n8999), .I1(n4_adj_197));
    OR3 i6508 (.O(n9154), .I0(n16_adj_39), .I1(n9123), .I2(n14_adj_83));
    AND2 i6688 (.O(n9338), .I0(n5812), .I1(n4459));
    OR2 i6458 (.O(n9100), .I0(key_in_c_0), .I1(n5874));
    AND4 i6624 (.O(n9274), .I0(n9279), .I1(n20_adj_1), .I2(n31), .I3(n25));
    XOR2 i6577 (.O(n9227), .I0(flag_Data[1]), .I1(flag_Data[0]));
    AND2 i6631 (.O(n9281), .I0(n15_adj_45), .I1(n9241));
    OR2 i6648 (.O(n9298), .I0(n9297), .I1(n9296));
    OR2 i6732 (.O(n9382), .I0(n9381), .I1(n9380));
    OR2 i6585 (.O(n5826), .I0(n9234), .I1(n9233));
    AND2 i6685 (.O(n9335), .I0(n5812), .I1(n8388));
    AND2 i6682 (.O(n9332), .I0(n8386), .I1(led_int_Data0_3__N_388[1]));
    AND2 i6679 (.O(n9329), .I0(n8386), .I1(led_int_Data0_3__N_388[2]));
    AND6 i6568 (.O(n9219), .I0(timecnt[3]), .I1(n9188), .I2(timecnt[2]), 
         .I3(n9082), .I4(timecnt[1]), .I5(timecnt[13]));
    OR2 i6632 (.O(n9282), .I0(n9281), .I1(n9280));
    OR2 key_in_3__I_0_244_i15 (.O(n15_adj_108), .I0(n14), .I1(n11_adj_115));
    OR2 i6516 (.O(n9162), .I0(n9005), .I1(n9146));
    AND2 i6676 (.O(n9326), .I0(n8386), .I1(led_int_Data0_3__N_388[3]));
    OR2 i6518 (.O(n9164), .I0(n22_adj_112), .I1(n9_adj_47));
    OR2 i1_adj_52 (.O(n38), .I0(n6141), .I1(n6225));
    AND2 i6650 (.O(n9300), .I0(n1464), .I1(n8680));
    OR2 i2_adj_53 (.O(n5841), .I0(n4_adj_48), .I1(flag_Data[0]));
    XOR2 i1113 (.O(led_int_Data0_3__N_388[1]), .I0(n3206), .I1(int_Data[1]));
    OR2 i2_adj_54 (.O(n4572), .I0(n9113), .I1(n783));
    OR2 key_in_3__I_0_245_i15 (.O(n15_adj_102), .I0(n14_adj_114), .I1(n11_adj_46));
    AND2 i3248 (.O(n5829), .I0(n15_adj_119), .I1(n15_adj_102));
    AND2 i1_adj_55 (.O(n8976), .I0(n6038), .I1(int_Data[2]));
    AND2 i6734 (.O(n9384), .I0(n1299), .I1(n535));
    OR2 i6522 (.O(n9168), .I0(n22_adj_19), .I1(n16));
    OR2 i1_adj_56 (.O(n8948), .I0(n8336), .I1(n104_adj_32));
    OR2 i6735 (.O(n9385), .I0(n9384), .I1(n9383));
    AND2 i5330 (.O(n7953), .I0(n7946), .I1(int_Data0[5]));
    XOR2 i2_adj_57 (.O(n8388), .I0(n4), .I1(n6_adj_23));
    OR3 i2_adj_58 (.O(n22_adj_130), .I0(n25), .I1(n18_adj_153), .I2(n21_adj_69));
    AND2 i1_adj_59 (.O(n8326), .I0(n8976), .I1(int_Data[5]));
    AND2 i2_adj_60 (.O(n84), .I0(n6_adj_24), .I1(n90_adj_118));
    OR2 i6651 (.O(n9301), .I0(n9300), .I1(n9299));
    XOR2 i1_adj_61 (.O(n9027), .I0(int_Data0[2]), .I1(int_Data1[2]));
    XOR2 i1_adj_62 (.O(n9028), .I0(n9027), .I1(n4_adj_168));
    AND2 i6530 (.O(n9178), .I0(n9123), .I1(n22_adj_42));
    AND4 i6532 (.O(n9180), .I0(n15_adj_106), .I1(n8982), .I2(n5916), 
         .I3(n15_adj_108));
    OR2 i6543 (.O(n9192), .I0(n9102), .I1(n9178));
    DFFCR int_Data__i1 (.Q(led_int_Data0_3__N_388[0]), .D(n9267), .CLK(time10ms), 
          .CE(n4698), .R(reset_c));   // calculate.v(55[13] 193[16])
    DFFR led_int_Data1_i4 (.Q(led_int_Data1_c_3), .D(led_int_Data1_3__N_63[3]), 
         .CLK(clk_c), .R(reset_c));   // calculate.v(204[13] 242[16])
    AND2 i6737 (.O(n9387), .I0(n1298), .I1(n525));
    AND2 i2_adj_63 (.O(n28_adj_151), .I0(n4_adj_85), .I1(n34_adj_144));
    XOR2 i2_adj_64 (.O(led_int_Data0_3__N_388[2]), .I0(n4_adj_198), .I1(n3504));
    AND2 i2_adj_65 (.O(n8335), .I0(n91_adj_31), .I1(n29_adj_29));
    OR2 i1_adj_66 (.O(n5999), .I0(n9022), .I1(n16_adj_39));
    IBUF key_in_pad_0 (.O(key_in_c_0), .I0(key_in[0]));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(186[8:12])
    IBUF key_in_pad_1 (.O(key_in_c_1), .I0(key_in[1]));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(186[8:12])
    IBUF key_in_pad_2 (.O(key_in_c_2), .I0(key_in[2]));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(186[8:12])
    XOR2 i1_adj_67 (.O(n8429), .I0(n9027), .I1(n4_adj_129));
    OR2 i5378 (.O(n8_adj_172), .I0(n8001), .I1(n8005));
    AND2 i6594 (.O(led_int_Data2_3__N_67[0]), .I0(n9243), .I1(n9242));
    AND2 i2_adj_68 (.O(n3187), .I0(n6_adj_86), .I1(n68_adj_145));
    IBUF key_in_pad_3 (.O(key_in_c_3), .I0(key_in[3]));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(186[8:12])
    IBUF reset_pad (.O(reset_c), .I0(reset));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(186[8:12])
    IBUF clk_pad (.O(clk_c), .I0(clk));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(186[8:12])
    OBUF key_out_pad_0 (.O(key_out[0]), .I0(key_out_c_0));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF key_out_pad_1 (.O(key_out[1]), .I0(key_out_c_1));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF key_out_pad_2 (.O(key_out[2]), .I0(key_out_c_2));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF key_out_pad_3 (.O(key_out[3]), .I0(key_out_c_3));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF led_int_Data2_pad_0 (.O(led_int_Data2[0]), .I0(led_int_Data2_c_0));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    AND2 i1_adj_69 (.O(n1_adj_196), .I0(n31), .I1(n84));
    OR2 i1_adj_70 (.O(n4_adj_197), .I0(n4546), .I1(n1_adj_196));
    OBUF led_int_Data2_pad_1 (.O(led_int_Data2[1]), .I0(led_int_Data2_c_3));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    AND3 i6764 (.O(n9414), .I0(key_in_c_2), .I1(n9413), .I2(n6_adj_187));
    OBUF led_int_Data2_pad_2 (.O(led_int_Data2[2]), .I0(n929));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OR2 i2_adj_71 (.O(n4588), .I0(n8341), .I1(n4587));
    AND2 i6619 (.O(n9269), .I0(key_out_c_3), .I1(n4_adj_97));
    OBUF led_int_Data2_pad_3 (.O(led_int_Data2[3]), .I0(led_int_Data2_c_3));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF led_int_Data1_pad_0 (.O(led_int_Data1[0]), .I0(led_int_Data1_c_0));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF led_int_Data1_pad_1 (.O(led_int_Data1[1]), .I0(led_int_Data1_c_1));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF led_int_Data1_pad_2 (.O(led_int_Data1[2]), .I0(led_int_Data1_c_2));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF led_int_Data1_pad_3 (.O(led_int_Data1[3]), .I0(led_int_Data1_c_3));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OR2 i1_adj_72 (.O(n9007), .I0(n9005), .I1(n22));
    AND2 i6653 (.O(n9303), .I0(n1464), .I1(n8642));
    AND4 i6549 (.O(n9198), .I0(n8979), .I1(n15_adj_6), .I2(n5883), .I3(n5820));
    DFFR led_int_Data1_i3 (.Q(led_int_Data1_c_2), .D(led_int_Data1_3__N_63[2]), 
         .CLK(clk_c), .R(reset_c));   // calculate.v(204[13] 242[16])
    DFFR led_int_Data1_i2 (.Q(led_int_Data1_c_1), .D(led_int_Data1_3__N_63[1]), 
         .CLK(clk_c), .R(reset_c));   // calculate.v(204[13] 242[16])
    DFFCR int_Data0_i0_i7 (.Q(int_Data0[7]), .D(n8343), .CLK(time10ms), 
          .CE(n4679), .R(reset_c));   // calculate.v(55[13] 193[16])
    DFFCR int_Data0_i0_i6 (.Q(int_Data0[6]), .D(n8352), .CLK(time10ms), 
          .CE(n4679), .R(reset_c));   // calculate.v(55[13] 193[16])
    OBUF led_int_Data0_pad_0 (.O(led_int_Data0[0]), .I0(led_int_Data0_c_0));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF led_int_Data0_pad_1 (.O(led_int_Data0[1]), .I0(led_int_Data0_c_1));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF led_int_Data0_pad_2 (.O(led_int_Data0[2]), .I0(led_int_Data0_c_2));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OR2 i6551 (.O(n9200), .I0(n9005), .I1(n9140));
    OBUF led_int_Data0_pad_3 (.O(led_int_Data0[3]), .I0(led_int_Data0_c_3));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OR2 i1_adj_73 (.O(n5835), .I0(n9005), .I1(n22_adj_130));
    DFFCR int_Data0_i0_i5 (.Q(int_Data0[5]), .D(n8349), .CLK(time10ms), 
          .CE(n4679), .R(reset_c));   // calculate.v(55[13] 193[16])
    DFFCR int_Data0_i0_i4 (.Q(int_Data0[4]), .D(n8348), .CLK(time10ms), 
          .CE(n4679), .R(reset_c));   // calculate.v(55[13] 193[16])
    DFFCR int_Data0_i0_i3 (.Q(int_Data0[3]), .D(n17_adj_35), .CLK(time10ms), 
          .CE(n4679), .R(reset_c));   // calculate.v(55[13] 193[16])
    OBUF PointTime_pad (.O(PointTime), .I0(PointTime_c));   // E:/Bin/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    DFFCR int_Data0_i0_i2 (.Q(int_Data0[2]), .D(n4588), .CLK(time10ms), 
          .CE(n4679), .R(reset_c));   // calculate.v(55[13] 193[16])
    DFFCR int_Data0_i0_i1 (.Q(int_Data0[1]), .D(n13_adj_41), .CLK(time10ms), 
          .CE(n4679), .R(reset_c));   // calculate.v(55[13] 193[16])
    DFFCS led_int_Data2_i4 (.Q(led_int_Data2_c_3), .D(led_int_Data2_3__N_67[3]), 
          .CLK(time10ms), .CE(n9282), .S(reset_c));   // calculate.v(55[13] 193[16])
    AND2 i6634 (.O(n9284), .I0(flag_Data[0]), .I1(n74_adj_52));
    DFFC key_out_i0_i4 (.Q(key_out_c_3), .D(scanvalue[3]), .CLK(time10ms), 
         .CE(reset_c));   // calculate.v(55[13] 193[16])
    OR4 i3_adj_74 (.O(n8354), .I0(n4558), .I1(flag_Cal[1]), .I2(n4_adj_97), 
        .I3(n78_adj_33));
    OR2 i3642 (.O(n6026), .I0(flag_Data[0]), .I1(n16));
    DFFC key_out_i0_i3 (.Q(key_out_c_2), .D(scanvalue[2]), .CLK(time10ms), 
         .CE(reset_c));   // calculate.v(55[13] 193[16])
    DFFC key_out_i0_i2 (.Q(key_out_c_1), .D(scanvalue[1]), .CLK(time10ms), 
         .CE(reset_c));   // calculate.v(55[13] 193[16])
    DFFCR flag_Data_i1 (.Q(flag_Data[1]), .D(n5795), .CLK(time10ms), .CE(n4712), 
          .R(reset_c));   // calculate.v(55[13] 193[16])
    AND2 i6554 (.O(n9203), .I0(n796), .I1(n9202));
    OR2 i1_adj_75 (.O(n4684), .I0(led_int_Data2_3__N_109), .I1(n9065));
    OR2 i6555 (.O(n4355), .I0(n770), .I1(n9203));
    OR2 i6590 (.O(n5856), .I0(n9239), .I1(n9238));
    AND2 i6561 (.O(n9211), .I0(n9200), .I1(n15_adj_73));
    AND3 i2_adj_76 (.O(n8452), .I0(n5_adj_93), .I1(n28), .I2(n31));
    AND2 i1115 (.O(n3504), .I0(n3206), .I1(int_Data[1]));
    INV i5827 (.O(n8467), .I0(n10_adj_18));
    AND2 i6765 (.O(n9415), .I0(n4548), .I1(n3_adj_186));
    AND4 i6565 (.O(n9217), .I0(n9164), .I1(n9148), .I2(n9168), .I3(n4_adj_48));
    OR4 i3_adj_77 (.O(n1_adj_185), .I0(key_in_c_0), .I1(key_out_c_0), 
        .I2(n4391), .I3(n7_adj_89));
    AND2 i1124 (.O(n3513), .I0(n3504), .I1(n3205));
    AND6 i6574 (.O(n5869), .I0(n9152), .I1(n9218), .I2(n9162), .I3(n9150), 
         .I4(n9154), .I5(n6181));
    OR2 i1125 (.O(n4148), .I0(n3504), .I1(n3205));
    INV i5828 (.O(n8468), .I0(n4492));
    OR2 i2_adj_78 (.O(n14_adj_107), .I0(n4_adj_195), .I1(n13));
    AND2 i1_adj_79 (.O(n4686), .I0(n9012), .I1(n4684));
    INV i5840 (.O(n8480), .I0(n14_adj_116));
    OR2 i6635 (.O(n9285), .I0(n9284), .I1(n9283));
    OR2 i6567 (.O(n9218), .I0(n9217), .I1(flag_Data[0]));
    OR2 i6597 (.O(n1480), .I0(n9246), .I1(n8305));
    DFFCR int_Data1_i0_i3 (.Q(int_Data1[3]), .D(n4651), .CLK(time10ms), 
          .CE(n4679), .R(reset_c));   // calculate.v(55[13] 193[16])
    AND2 i6599 (.O(n4698), .I0(n9248), .I1(n85));
    AND2 i1_adj_80 (.O(n35), .I0(n9013), .I1(key_in_c_2));
    OR2 i6617 (.O(n9267), .I0(n9266), .I1(n9265));
    AND2 i6621 (.O(n9271), .I0(n3842), .I1(led_int_Data2_3__N_111[1]));
    OR2 i6654 (.O(n9304), .I0(n9303), .I1(n9302));
    OR2 i1_adj_81 (.O(n15_adj_194), .I0(n4567), .I1(n1_adj_192));
    AND2 i6602 (.O(n8364), .I0(n9251), .I1(n9250));
    AND3 i3_adj_82 (.O(n8305), .I0(n9319), .I1(n82_adj_51), .I2(n5_adj_110));
    AND2 i1_adj_83 (.O(n41), .I0(n9_adj_47), .I1(key_out_c_2));
    AND3 i6656 (.O(n9306), .I0(n6_adj_99), .I1(key_in_c_1), .I2(n4_adj_70));
    AND2 i6605 (.O(n17_adj_35), .I0(n9254), .I1(n9253));
    OR3 i1_adj_84 (.O(n8953), .I0(n6042), .I1(n43), .I2(key_in_c_0));
    OR2 key_in_3__I_0_246_i15 (.O(n15_adj_87), .I0(n14_adj_74), .I1(n11_adj_7));
    AND2 i2_adj_85 (.O(n82), .I0(n4_adj_100), .I1(n87_adj_109));
    AND2 i6637 (.O(n9287), .I0(n9286), .I1(n540));
    OR2 i6608 (.O(led_int_Data2_3__N_67[3]), .I0(n9257), .I1(n9256));
    OR3 i1_adj_86 (.O(n8955), .I0(n9_adj_160), .I1(n1_adj_179), .I2(n1323));
    OR2 key_in_3__I_0_237_i15 (.O(n15_adj_11), .I0(n14_adj_107), .I1(n11_adj_7));
    AND2 i3243 (.O(n96), .I0(n29), .I1(n79_adj_127));
    AND2 i6618 (.O(n9268), .I0(n32_adj_30), .I1(n20));
    AND2 i6638 (.O(n9288), .I0(n9118), .I1(n7911));
    OR2 i2_adj_87 (.O(n4520), .I0(n4_adj_157), .I1(led_int_Data1_3__N_385));
    OR2 i1_adj_88 (.O(n5839), .I0(n9022), .I1(n16));
    XOR2 i5463 (.O(n73_adj_105), .I0(n8085), .I1(timecnt[7]));
    AND2 i6611 (.O(n4679), .I0(n9260), .I1(n9259));
    OR2 i3505 (.O(n6099), .I0(n5955), .I1(n537));
    AND2 i5379 (.O(n8005), .I0(n8004), .I1(int_Data0[3]));
    OR2 i1_adj_89 (.O(n9013), .I0(key_in_c_1), .I1(key_in_c_0));
    AND3 i2_adj_90 (.O(n8352), .I0(n9040), .I1(int_Data0[6]), .I2(flag_Data[1]));
    OR3 i1_adj_91 (.O(n8959), .I0(n16_adj_193), .I1(n757), .I2(n770));
    AND2 i6614 (.O(n19_adj_188), .I0(n9263), .I1(n9262));
    OR2 i6657 (.O(n9307), .I0(n9306), .I1(n9305));
    AND3 i6659 (.O(n9309), .I0(n4549), .I1(key_in_c_0), .I2(n87_adj_109));
    AND2 i3446 (.O(n6038), .I0(int_Data[3]), .I1(int_Data[4]));
    OR2 i6639 (.O(n9289), .I0(n9288), .I1(n9287));
    AND2 i5642 (.O(n8281), .I0(n8280), .I1(n3722));
    AND3 i1_adj_92 (.O(n8961), .I0(n8473), .I1(int_Data1_7__N_351[3]), 
         .I2(n8444));
    AND4 i1_adj_93 (.O(n8963), .I0(n6214), .I1(n15_adj_40), .I2(n15_adj_113), 
         .I3(n15_adj_11));
    AND3 i2_adj_94 (.O(n8341), .I0(n9045), .I1(int_Data0[2]), .I2(flag_Data[1]));
    INV i46 (.O(n6581), .I0(n9004));
    OR2 i3450 (.O(n6042), .I0(key_in_c_3), .I1(key_out_c_3));
    AND3 i1_adj_95 (.O(n8964), .I0(n8988), .I1(n8457), .I2(n8_adj_21));
    OR2 i6660 (.O(n9310), .I0(n9309), .I1(n9308));
    AND2 i1_adj_96 (.O(n4712), .I0(n4680), .I1(n8598));
    OR2 i1_adj_97 (.O(n28), .I0(key_out_c_1), .I1(n29_adj_29));
    AND3 i6662 (.O(n9312), .I0(n4543), .I1(key_in_c_3), .I2(key_out_c_2));
    AND3 i2_adj_98 (.O(n8302), .I0(n15_adj_102), .I1(n97), .I2(n5953));
    AND3 i2_adj_99 (.O(n4546), .I0(n31), .I1(n87_adj_109), .I2(n4_adj_100));
    AND2 i3242 (.O(n95), .I0(n29), .I1(n78));
    AND2 i1_adj_100 (.O(n9065), .I0(n85), .I1(n9064));
    OR2 key_in_3__I_0_248_i14 (.O(n14_adj_74), .I0(n16_adj_91), .I1(n9013));
    OR2 i6766 (.O(n9416), .I0(n9415), .I1(n9414));
    AND2 i1046 (.O(n3435), .I0(n4_adj_14), .I1(n1556));
    OR2 i6663 (.O(n99), .I0(n9312), .I1(n9311));
    AND2 i6496 (.O(n9142), .I0(n50), .I1(n49_adj_150));
    OR2 i1048 (.O(n6_adj_23), .I0(n3435), .I1(n8345));
    AND2 i6767 (.O(n9417), .I0(n9250), .I1(n9416));
    AND4 i1_adj_101 (.O(n4_adj_65), .I0(n15_adj_8), .I1(n5926), .I2(n94), 
         .I3(n15_adj_133));
    AND3 i2_adj_102 (.O(n8318), .I0(n9310), .I1(n25), .I2(n10));
    AND2 i3288 (.O(n1466), .I0(n5869), .I1(n9376));
    AND2 i1013 (.O(n14_adj_116), .I0(int_Data[6]), .I1(n4567));
    AND2 i3239 (.O(n6101), .I0(n11_adj_115), .I1(n11_adj_10));
    AND2 i2_adj_103 (.O(n109), .I0(n4_adj_70), .I1(n108));
    AND3 i6665 (.O(n9315), .I0(n6_adj_86), .I1(key_in_c_0), .I2(n97_adj_28));
    AND2 i3454 (.O(n6191), .I0(n17), .I1(n6026));
    AND2 i6622 (.O(n9272), .I0(flag_Data[1]), .I1(int_Data0[1]));
    OR2 i6666 (.O(n9316), .I0(n9315), .I1(n9314));
    OR3 i2_adj_104 (.O(n6214), .I0(n10_adj_121), .I1(n14), .I2(n9102));
    OR2 i3235 (.O(led_int_Data1_3__N_63[0]), .I0(led_int_Data1_3__N_385), 
        .I1(led_int_Data1_3__N_381[0]));
    OR2 key_in_3__I_0_249_i15 (.O(n15_adj_53), .I0(n14_adj_107), .I1(n11_adj_46));
    OR2 i6738 (.O(n9388), .I0(n9387), .I1(n9386));
    AND2 i1_adj_105 (.O(n25_adj_190), .I0(n24_adj_189), .I1(n9063));
    AND2 i3234 (.O(led_int_Data1_3__N_381[0]), .I0(n1524), .I1(n874));
    OR2 i1_adj_106 (.O(n9012), .I0(n9010), .I1(flag_Cal[1]));
    AND2 i3370 (.O(n6189), .I0(n6141), .I1(n14_adj_114));
    OR2 i1_adj_107 (.O(n9008), .I0(n9005), .I1(n22_adj_75));
    OR2 i1_adj_108 (.O(n9010), .I0(flag_Cal[0]), .I1(n15_adj_45));
    XOR2 i1_adj_109 (.O(n9030), .I0(int_Data0[3]), .I1(int_Data1[3]));
    AND2 i6526 (.O(n9172), .I0(timecnt[10]), .I1(timecnt[5]));
    INV i6578 (.O(n1701), .I0(n9227));
    INV i6580 (.O(n9230), .I0(n4_adj_124));
    OR2 i3233 (.O(n874), .I0(n744), .I1(n864));
    AND2 i6673 (.O(n9323), .I0(n3842), .I1(n19_adj_37));
    AND2 i6539 (.O(n9188), .I0(n9172), .I1(timecnt[8]));
    INV i6589 (.O(n9239), .I0(n15_adj_87));
    AND2 i1_adj_110 (.O(n8978), .I0(n8976), .I1(int_Data[1]));
    INV i6553 (.O(n9202), .I0(n783));
    INV i14 (.O(n8744), .I0(n8959));
    INV i6595 (.O(n9245), .I0(time10ms));
    OR2 key_in_3__I_0_250_i15 (.O(n15_adj_44), .I0(n14), .I1(n11_adj_46));
    INV i6596 (.O(n9246), .I0(n15_adj_45));
    OR3 i2_adj_111 (.O(n5843), .I0(n16_adj_39), .I1(n22_adj_146), .I2(flag_Data[0]));
    INV i4_adj_112 (.O(n8477), .I0(int_Data[7]));
    INV i6598 (.O(n9248), .I0(n8948));
    OR2 equal_413_i19 (.O(n19_adj_25), .I0(n18), .I1(n25));
    INV i1_adj_113 (.O(n1_adj_192), .I0(n4564));
    AND2 i6740 (.O(n9390), .I0(n1299), .I1(n536));
    INV i6600 (.O(n9250), .I0(n3187));
    INV i6601 (.O(n9251), .I0(n4_adj_61));
    AND3 i6668 (.O(n9318), .I0(n5_adj_93), .I1(key_in_c_3), .I2(n92_adj_147));
    INV i6603 (.O(n9253), .I0(n29_adj_34));
    OR2 i6669 (.O(n9319), .I0(n9318), .I1(n9317));
    OR2 i3230 (.O(n854), .I0(n770), .I1(n796));
    AND2 i6494 (.O(n9140), .I0(n9068), .I1(n22_adj_75));
    OR2 i1_adj_114 (.O(n8712), .I0(n10_adj_9), .I1(n7));
    OR2 i3507 (.O(n5820), .I0(n6101), .I1(n14_adj_107));
    INV i6604 (.O(n9254), .I0(n9325));
    INV i6606 (.O(n9256), .I0(flag_Data[0]));
    INV i6607 (.O(n9257), .I0(n5795));
    INV i6609 (.O(n9259), .I0(n64));
    AND2 i6768 (.O(n9418), .I0(n3187), .I1(n1_adj_185));
    AND3 i2_adj_115 (.O(n8340), .I0(n9051), .I1(int_Data1[1]), .I2(n5887));
    INV i6610 (.O(n9260), .I0(n67_adj_78));
    INV i6612 (.O(n9262), .I0(n25_adj_190));
    INV i6575 (.O(n1464), .I0(n5869));
    INV i6613 (.O(n9263), .I0(n9419));
    INV i6497 (.O(n4_adj_135), .I0(n9142));
    AND3 i1_adj_116 (.O(n10_adj_9), .I0(flag_Data[1]), .I1(n9), .I2(int_Data0[0]));
    AND2 i2_adj_117 (.O(n757), .I0(n4_adj_2), .I1(n8458));
    AND2 i2_adj_118 (.O(n731), .I0(n4_adj_184), .I1(n8468));
    INV i6493 (.O(n9), .I0(n9138));
    INV i6491 (.O(n6_adj_95), .I0(n9136));
    VCC i6576 (.X(pwr));
    OR2 i3228 (.O(n3206), .I0(led_int_Data1_3__N_385), .I1(n1524));
    AND3 i2_adj_119 (.O(n8339), .I0(n9060), .I1(int_Data1[2]), .I2(n5887));
    OR3 i1_adj_120 (.O(n8598), .I0(n9321), .I1(n9320), .I2(n1207));
    XOR2 i5491 (.O(n69_adj_123), .I0(n8113), .I1(timecnt[11]));
    XOR2 i1_adj_121 (.O(n4_adj_141), .I0(n8146), .I1(n34));
    XOR2 i5498 (.O(n68_adj_103), .I0(n8120), .I1(timecnt[12]));
    XOR2 i1_adj_122 (.O(n4_adj_149), .I0(n8_adj_62), .I1(n3722));
    AND2 i1_adj_123 (.O(n7), .I0(n6_adj_95), .I1(int_Data0_7__N_183[0]));
    XOR2 i1_adj_124 (.O(n4_adj_158), .I0(n5797), .I1(int_Data[2]));
    OR2 i6741 (.O(n9391), .I0(n9390), .I1(n9389));
    AND4 i1_adj_125 (.O(n9_adj_22), .I0(n5837), .I1(n5839), .I2(n5841), 
         .I3(n5835));
    XOR2 i5470 (.O(n72_adj_104), .I0(n8092), .I1(timecnt[8]));
    XOR2 i1_adj_126 (.O(n4_adj_161), .I0(n8_adj_175), .I1(n3757));
    XOR2 i1_adj_127 (.O(n4_adj_162), .I0(n8241), .I1(n3725));
    AND2 i3291 (.O(n1467), .I0(n5869), .I1(n9382));
    AND2 i5587 (.O(n8220), .I0(n8219), .I1(n3758));
    XOR2 i1_adj_128 (.O(n4_adj_166), .I0(n4_adj_76), .I1(n3724));
    INV i6557 (.O(n9045), .I0(n9205));
    XOR2 i1_adj_129 (.O(n4_adj_177), .I0(n6_adj_67), .I1(n3723));
    XOR2 i1_adj_130 (.O(n4_adj_178), .I0(n6_adj_165), .I1(n82_adj_60));
    OR2 i6769 (.O(n9419), .I0(n9418), .I1(n9417));
    INV i6484 (.O(n8996), .I0(n9128));
    OR2 i2_adj_131 (.O(n11_adj_46), .I0(n4_adj_97), .I1(n32_adj_30));
    INV i6480 (.O(n9060), .I0(n9124));
    INV i1_adj_132 (.O(n1_adj_179), .I0(n5839));
    XOR2 i5505 (.O(n67_adj_59), .I0(n8127), .I1(timecnt[13]));
    OR3 i2_adj_133 (.O(n9021), .I0(n8971), .I1(n3_adj_84), .I2(n9019));
    XOR2 i1_adj_134 (.O(n9031), .I0(n9030), .I1(n6_adj_164));
    INV i19 (.O(n6_adj_24), .I0(n9_adj_47));
    INV i20 (.O(led_int_Data2_3__N_111[1]), .I0(flag_Data[0]));
    INV i5800 (.O(n539), .I0(n8439));
    AND3 i2_adj_135 (.O(n8336), .I0(n4_adj_70), .I1(n6_adj_98), .I2(n100));
    INV i3496 (.O(n6089), .I0(n4520));
    AND2 i3232 (.O(n864), .I0(n5812), .I1(n854));
    INV i24_adj_136 (.O(n8642), .I0(n9018));
    INV i6763 (.O(n9413), .I0(n4548));
    OR2 i1_adj_137 (.O(n15_adj_40), .I0(n3842), .I1(n4_adj_65));
    OR2 i1_adj_138 (.O(n4_adj_97), .I0(key_out_c_2), .I1(n9_adj_47));
    INV i5867 (.O(n1489), .I0(n8506));
    INV i1929 (.O(n1490), .I0(n4464));
    INV i5804 (.O(n8444), .I0(n11_adj_115));
    AND2 i6500 (.O(n9146), .I0(n22_adj_130), .I1(n22));
    INV i1936 (.O(n1485), .I0(n4471));
    AND2 i6743 (.O(n9393), .I0(n1298), .I1(n526));
    AND2 i3227 (.O(n92_adj_43), .I0(n29), .I1(n75_adj_63));
    INV i3660 (.O(n1512), .I0(n8386));
    AND2 i3226 (.O(n91), .I0(n29), .I1(n74));
    INV i1938 (.O(n1486), .I0(n4473));
    OR2 i2_adj_139 (.O(n8386), .I0(n3205), .I1(n744));
    OR2 key_in_3__I_0_i15 (.O(n15_adj_45), .I0(n14_adj_74), .I1(n11_adj_46));
    OR2 i3372 (.O(n5955), .I0(n5861), .I1(n538));
    AND3 i2_adj_140 (.O(n8317), .I0(n99), .I1(n20_adj_1), .I2(n10));
    OR2 i3374 (.O(n5957), .I0(int_Data[5]), .I1(int_Data[4]));
    AND2 i3225 (.O(n90), .I0(n29), .I1(n73_adj_105));
    AND2 i5466 (.O(n8092), .I0(n8085), .I1(timecnt[7]));
    AND3 i6671 (.O(n9321), .I0(n1_adj_156), .I1(n7_adj_89), .I2(flag_Data[1]));
    OR2 i5302 (.O(n4_adj_168), .I0(n7920), .I1(n7924));
    XOR2 i5328 (.O(n525), .I0(n7946), .I1(int_Data0[5]));
    AND2 i5592 (.O(n8225), .I0(n8_adj_175), .I1(n124));
    AND2 i5303 (.O(n7924), .I0(n7923), .I1(int_Data0[1]));
    OR2 i5593 (.O(n8228), .I0(n8_adj_175), .I1(n124));
    OR2 i5594 (.O(n10_adj_174), .I0(n8225), .I1(n8229));
    XOR2 i5512 (.O(n66_adj_92), .I0(n8134), .I1(timecnt[14]));
    XOR2 i5335 (.O(n524), .I0(n7953), .I1(int_Data0[6]));
    INV i6591 (.O(n9241), .I0(n24));
    INV i1940 (.O(n1487), .I0(n4475));
    INV i3461 (.O(n4543), .I0(n6052));
    INV i6473 (.O(n9048), .I0(n9116));
    OR2 key_in_3__I_0_242_i13 (.O(n13), .I0(key_in_c_3), .I1(key_in_c_2));
    AND2 i3224 (.O(n89), .I0(n29), .I1(n72_adj_104));
    AND2 i3223 (.O(n88), .I0(n29), .I1(n71));
    INV i3451 (.O(n4549), .I0(n6042));
    AND2 i3334 (.O(n9086), .I0(n4_adj_195), .I1(n4_adj_64));
    INV i5833 (.O(n8473), .I0(n6141));
    OR6 i6_adj_141 (.O(n29), .I0(timecnt[7]), .I1(timecnt[11]), .I2(n10_adj_101), 
        .I3(timecnt[6]), .I4(timecnt[9]), .I5(n8950));
    XOR2 i1_adj_142 (.O(n8425), .I0(n9030), .I1(n6_adj_171));
    INV i5802 (.O(n536), .I0(n8441));
    INV i6550 (.O(n9040), .I0(n9198));
    INV i6582 (.O(n9232), .I0(n5826));
    AND2 i3222 (.O(n87), .I0(n29), .I1(n70));
    OR2 i6502 (.O(n9148), .I0(n16_adj_39), .I1(n22_adj_42));
    OR2 i6744 (.O(n9394), .I0(n9393), .I1(n9392));
    INV i6583 (.O(n9233), .I0(n15_adj_44));
    XOR2 i5342 (.O(n523), .I0(n7960), .I1(int_Data0[7]));
    INV sub_115_inv_0_i2 (.O(n8), .I0(int_Data1[1]));
    OR2 i1002 (.O(n8_adj_21), .I0(int_Data[3]), .I1(n6_adj_117));
    AND2 i3221 (.O(n86), .I0(n29), .I1(n69_adj_123));
    AND2 i999 (.O(n12_adj_71), .I0(int_Data[5]), .I1(n10_adj_79));
    OR2 i998 (.O(n10_adj_79), .I0(int_Data[4]), .I1(int_Data[3]));
    AND2 i3220 (.O(n85_adj_143), .I0(n29), .I1(n68_adj_103));
    AND2 i5473 (.O(n8099), .I0(n8092), .I1(timecnt[8]));
    AND2 i5445 (.O(n8071), .I0(n8064), .I1(timecnt[4]));
    OR2 i5386 (.O(n10_adj_170), .I0(n8_adj_172), .I1(int_Data0[4]));
    AND2 i6746 (.O(n9396), .I0(n1299), .I1(n537));
    AND2 i3219 (.O(n84_adj_131), .I0(n29), .I1(n67_adj_59));
    AND2 i1_adj_143 (.O(n9080), .I0(n11_adj_7), .I1(n11_adj_46));
    AND2 i5520 (.O(n8146), .I0(n31_adj_50), .I1(n11_adj_155));
    AND2 i5595 (.O(n8229), .I0(n8228), .I1(n3757));
    OR2 i6747 (.O(n9397), .I0(n9396), .I1(n9395));
    AND2 i1_adj_144 (.O(n4548), .I0(n8999), .I1(n4546));
    INV sub_115_inv_0_i3 (.O(n7_adj_13), .I0(int_Data1[2]));
    INV sub_115_inv_0_i4 (.O(n6), .I0(int_Data1[3]));
    XOR2 i1_adj_145 (.O(n4_adj_198), .I0(int_Data[2]), .I1(n3205));
    INV i1348 (.O(n3830), .I0(n4067));
    XOR2 i1_adj_146 (.O(n4), .I0(n4355), .I1(int_Data[3]));
    INV i3_adj_147 (.O(n3_adj_84), .I0(n22_adj_130));
    INV i5858 (.O(n8498), .I0(n8978));
    XOR2 i5477 (.O(n71), .I0(n8099), .I1(timecnt[9]));
    OR2 i5530 (.O(n8158), .I0(n8146), .I1(n55_adj_134));
    INV i15 (.O(n15_adj_81), .I0(n4555));
    OR3 i2_adj_148 (.O(n22_adj_75), .I0(n32_adj_30), .I1(n4555), .I2(n31));
    AND2 i5529 (.O(n8155), .I0(n8146), .I1(n55_adj_134));
    AND3 i2_adj_149 (.O(n4_adj_68), .I0(n50), .I1(n4_adj_85), .I2(n34_adj_144));
    AND2 i6641 (.O(n9291), .I0(flag_Data[1]), .I1(int_Data0[0]));
    OR2 i5394 (.O(n12), .I0(n10_adj_170), .I1(int_Data0[5]));
    OR2 i5569 (.O(n8201), .I0(n8189), .I1(n52));
    AND2 i5360 (.O(n7983), .I0(n2), .I1(n8));
    AND2 i5308 (.O(n7929), .I0(n4_adj_168), .I1(int_Data1[2]));
    AND2 i6749 (.O(n9399), .I0(n1298), .I1(n9031));
    OR2 i5309 (.O(n7932), .I0(n4_adj_168), .I1(int_Data1[2]));
    OR2 i1_adj_150 (.O(n4609), .I0(n4608), .I1(n8313));
    OR2 i5531 (.O(n4_adj_163), .I0(n8155), .I1(n8159));
    AND2 i5532 (.O(n8159), .I0(n8158), .I1(n34));
    AND3 i2_adj_151 (.O(n8980), .I0(n5992), .I1(n6107), .I2(n8979));
    OR2 i5402 (.O(n14_adj_169), .I0(n12), .I1(int_Data0[6]));
    AND2 i5647 (.O(n8286), .I0(n10_adj_58), .I1(n145));
    OR2 i5310 (.O(n6_adj_164), .I0(n7929), .I1(n7933));
    OR2 i5648 (.O(n8289), .I0(n10_adj_58), .I1(n145));
    AND2 i5537 (.O(n8164), .I0(n4_adj_163), .I1(n79_adj_111));
    OR2 i5649 (.O(n12_adj_55), .I0(n8286), .I1(n8290));
    AND2 i5559 (.O(n8189), .I0(n28_adj_5), .I1(n8_adj_38));
    AND2 i990 (.O(n6_adj_137), .I0(int_Data[2]), .I1(int_Data[1]));
    OR2 i5538 (.O(n8167), .I0(n4_adj_163), .I1(n79_adj_111));
    AND2 i5459 (.O(n8085), .I0(n8078), .I1(timecnt[6]));
    INV i6466 (.O(n4_adj_96), .I0(n9108));
    INV i6464 (.O(n9054), .I0(n9106));
    INV i39 (.O(n9_adj_82), .I0(n7_adj_89));
    INV i43 (.O(n43), .I0(n100));
    INV i47 (.O(n47), .I0(n102));
    INV i6544 (.O(n79_adj_54), .I0(n9192));
    INV i5818 (.O(n8458), .I0(n4561));
    INV i6459 (.O(n5_adj_110), .I0(n9100));
    INV i6457 (.O(n9057), .I0(n9098));
    INV i6584 (.O(n9234), .I0(n15_adj_87));
    OR2 i5586 (.O(n8_adj_175), .I0(n8216), .I1(n8220));
    INV sub_115_inv_0_i1 (.O(n9_adj_26), .I0(int_Data1[0]));
    INV i5786 (.O(n537), .I0(n8425));
    INV i2119 (.O(n4680), .I0(n8360));
    INV i4_adj_152 (.O(n4_adj_36), .I0(int_Data0[3]));
    AND3 i2_adj_153 (.O(n8979), .I0(n6093), .I1(n15_adj_102), .I2(n6020));
    AND2 i986 (.O(n10_adj_18), .I0(int_Data[4]), .I1(n8_adj_15));
    OR2 i6504 (.O(n9150), .I0(n6191), .I1(n22_adj_146));
    OR2 i985 (.O(n8_adj_15), .I0(int_Data[3]), .I1(int_Data[2]));
    AND2 i5311 (.O(n7933), .I0(n7932), .I1(int_Data0[2]));
    AND2 i5568 (.O(n8198), .I0(n8189), .I1(n52));
    XOR2 i1_adj_154 (.O(n4_adj_176), .I0(n8189), .I1(n3760));
    AND2 i6581 (.O(led_int_Data1_3__N_63[3]), .I0(n9230), .I1(n9229));
    XOR2 i5289 (.O(n540), .I0(int_Data1[0]), .I1(int_Data0[0]));
    OR2 i5539 (.O(n6_adj_165), .I0(n8164), .I1(n8168));
    AND2 i5540 (.O(n8168), .I0(n8167), .I1(n58));
    OR2 i6750 (.O(n9400), .I0(n9399), .I1(n9398));
    AND2 i1_adj_155 (.O(n106_adj_80), .I0(n9307), .I1(n29_adj_29));
    AND2 i1_adj_156 (.O(n4554), .I0(n4_adj_94), .I1(n92_adj_147));
    XOR2 i5484 (.O(n70), .I0(n8106), .I1(timecnt[10]));
    OR2 i1_adj_157 (.O(n108), .I0(n8317), .I1(n8335));
    AND3 i1_adj_158 (.O(n8991), .I0(n15_adj_113), .I1(n15_adj_133), .I2(n15_adj_8));
    OR2 i1_adj_159 (.O(n4555), .I0(n21_adj_69), .I1(key_out_c_2));
    OR2 i5616 (.O(n8253), .I0(n8241), .I1(n49));
    AND2 i6752 (.O(n9402), .I0(n1299), .I1(n538));
    OR3 i2_adj_160 (.O(n3_adj_186), .I0(n7_adj_89), .I1(n20_adj_1), .I2(key_in_c_2));
    AND2 i5606 (.O(n8241), .I0(n25_adj_159), .I1(n5));
    AND2 i5615 (.O(n8250), .I0(n8241), .I1(n49));
    XOR2 i1_adj_161 (.O(time10ms_N_397), .I0(n29), .I1(n9245));
    AND2 i5452 (.O(n8078), .I0(n8071), .I1(timecnt[5]));
    OR2 i5410 (.O(n531), .I0(n14_adj_169), .I1(int_Data0[7]));
    OR2 equal_415_i18 (.O(n18), .I0(key_in_c_0), .I1(key_out_c_3));
    AND2 i5584 (.O(n8216), .I0(n6_adj_182), .I1(n100_adj_128));
    AND2 i6615 (.O(n9265), .I0(n5869), .I1(n9289));
    OR2 i5301 (.O(n7923), .I0(n7911), .I1(int_Data1[1]));
    OR2 i6753 (.O(n9403), .I0(n9402), .I1(n9401));
    OR2 i5354 (.O(n2), .I0(n9_adj_26), .I1(int_Data0[0]));
    OR2 i5361 (.O(n7986), .I0(n2), .I1(n8));
    OR2 i1_adj_162 (.O(n111), .I0(n106_adj_80), .I1(n8318));
    OR2 i1_adj_163 (.O(n85), .I0(n112), .I1(n109));
    AND3 i2_adj_164 (.O(n8349), .I0(n4787), .I1(int_Data0[5]), .I2(flag_Data[1]));
    AND2 i6460 (.O(n9102), .I0(n16_adj_39), .I1(n16));
    OR2 i5362 (.O(n4_adj_129), .I0(n7983), .I1(n7987));
    AND2 i1_adj_165 (.O(n112), .I0(n111), .I1(n9_adj_27));
    AND2 i3512 (.O(n6107), .I0(n5850), .I1(n15_adj_106));
    OR6 i6_adj_166 (.O(n8360), .I0(n9269), .I1(n32), .I2(n10_adj_180), 
        .I3(n8_adj_181), .I4(n9268), .I5(n26));
    AND2 i978 (.O(n8_adj_126), .I0(int_Data[3]), .I1(n6_adj_117));
    AND2 i5363 (.O(n7987), .I0(n7986), .I1(int_Data0[1]));
    AND2 i6441 (.O(n9082), .I0(timecnt[12]), .I1(timecnt[14]));
    OR2 i3_adj_167 (.O(n10_adj_101), .I0(n80), .I1(timecnt[4]));
    OR2 i1_adj_168 (.O(n8_adj_181), .I0(n15), .I1(n41));
    XOR2 i1_adj_169 (.O(n8_adj_77), .I0(n12_adj_55), .I1(n106));
    INV i6451 (.O(n9063), .I0(n9092));
    INV i6586 (.O(n9236), .I0(n8963));
    INV i6424 (.O(n9064), .I0(n28_adj_122));
    XOR2 i1_adj_170 (.O(n4_adj_90), .I0(n10_adj_58), .I1(n3721));
    INV i1188 (.O(n29_adj_29), .I0(key_in_c_3));
    XOR2 i1_adj_171 (.O(n4_adj_17), .I0(n4_adj_163), .I1(n58));
    INV i1_adj_172 (.O(n1_adj_156), .I0(n79));
    XOR2 i1_adj_173 (.O(n4_adj_152), .I0(n4_adj_183), .I1(n3759));
    INV i6592 (.O(n9242), .I0(n531));
    INV i3590 (.O(n4607), .I0(n8993));
    INV i1182 (.O(n32_adj_30), .I0(key_out_c_3));
    INV i3340 (.O(n1208), .I0(n5921));
    INV i16 (.O(n8680), .I0(n9017));
    INV key_in_3__I_0_i16 (.O(led_int_Data2_3__N_109), .I0(n15_adj_45));
    INV i3580 (.O(n1305), .I0(n6181));
    INV i5790 (.O(n538), .I0(n8429));
    OR2 i6506 (.O(n9152), .I0(n22_adj_19), .I1(n17));
    INV i5788 (.O(n1491), .I0(n8427));
    INV equal_404_i20 (.O(n1298), .I0(n8354));
    INV i6569 (.O(n8950), .I0(n9219));
    INV equal_405_i22 (.O(n1299), .I0(n4491));
    INV i5794 (.O(n533), .I0(n8433));
    INV i1134 (.O(n31), .I0(key_in_c_0));
    INV i1_adj_174 (.O(n1), .I0(flag_Cal[1]));
    INV i5817 (.O(n8457), .I0(n8326));
    AND2 i5545 (.O(n8173), .I0(n6_adj_165), .I1(n103));
    AND2 i1_adj_175 (.O(n115), .I0(n104), .I1(n20_adj_1));
    XOR2 i148 (.O(n90_adj_118), .I0(key_out_c_3), .I1(key_out_c_2));
    AND2 i1_adj_176 (.O(n8988), .I0(int_Data[4]), .I1(int_Data[5]));
    AND3 i2_adj_177 (.O(n796), .I0(n9054), .I1(n14_adj_116), .I2(n8477));
    INV equal_406_i22 (.O(n1300), .I0(n4490));
    OR2 i5585 (.O(n8219), .I0(n6_adj_182), .I1(n100_adj_128));
    AND2 i5650 (.O(n8290), .I0(n8289), .I1(n3721));
    XOR2 i146 (.O(n87_adj_109), .I0(key_out_c_1), .I1(key_out_c_0));
    OR2 i2_adj_178 (.O(n14_adj_114), .I0(n4_adj_64), .I1(n13));
    AND2 i5300 (.O(n7920), .I0(n7911), .I1(int_Data1[1]));
    AND2 i5480 (.O(n8106), .I0(n8099), .I1(timecnt[9]));
    OR2 i1_adj_179 (.O(n8504), .I0(n8_adj_126), .I1(int_Data[4]));
    OR2 i1_adj_180 (.O(n4_adj_61), .I0(n4548), .I1(key_in_c_2));
    AND2 i6674 (.O(n9324), .I0(flag_Data[1]), .I1(n4_adj_36));
    INV i3748 (.O(n4789), .I0(n8980));
    OR2 i3_adj_181 (.O(n10_adj_180), .I0(n8452), .I1(n35));
    XOR2 i147 (.O(n104), .I0(key_in_c_2), .I1(key_in_c_1));
    OR3 i2_adj_182 (.O(n4558), .I0(n16_adj_91), .I1(n32_adj_30), .I2(n9013));
    XOR2 i2_adj_183 (.O(n3757), .I0(n4_adj_178), .I1(n103));
    XOR2 i1_adj_184 (.O(n9033), .I0(int_Data0[1]), .I1(int_Data1[1]));
    OR2 i6642 (.O(int_Data0_7__N_183[0]), .I0(n9291), .I1(n9290));
    AND2 i6463 (.O(n9106), .I0(int_Data[6]), .I1(n5957));
    OR2 i3460 (.O(n6052), .I0(key_in_c_2), .I1(key_out_c_1));
    XOR2 i1_adj_185 (.O(n8439), .I0(n9033), .I1(n2));
    OR3 i2_adj_186 (.O(n19_adj_37), .I0(n11_adj_115), .I1(flag_Data[0]), 
        .I2(n6141));
    AND2 i6670 (.O(n9320), .I0(n9_adj_82), .I1(n1208));
    AND3 i2_adj_187 (.O(n783), .I0(n8480), .I1(n4564), .I2(n8477));
    AND4 i2_adj_188 (.O(n29_adj_34), .I0(n5829), .I1(n38), .I2(n5916), 
         .I3(n6020));
    INV i3311 (.O(n4_adj_70), .I0(n18));
    INV i12 (.O(n12_adj_138), .I0(n108));
    XOR2 i1_adj_189 (.O(n8433), .I0(n14_adj_169), .I1(int_Data0[7]));
    INV i5796 (.O(n534), .I0(n8435));
    OR2 i1_adj_190 (.O(n22_adj_42), .I0(n4555), .I1(n18_adj_153));
    XOR2 i2_adj_191 (.O(n3724), .I0(n4_adj_176), .I1(n52));
    OR2 equal_406_i18 (.O(n16_adj_91), .I0(n29_adj_29), .I1(key_in_c_2));
    AND2 i5487 (.O(n8113), .I0(n8106), .I1(timecnt[10]));
    XOR2 i2_adj_192 (.O(n3722), .I0(n4_adj_191), .I1(n100_adj_128));
    AND3 i6644 (.O(n9294), .I0(n6181), .I1(n1464), .I2(n8996));
    AND2 i5368 (.O(n7992), .I0(n4_adj_129), .I1(n7_adj_13));
    XOR2 i2_adj_193 (.O(n3723), .I0(n4_adj_152), .I1(n76));
    AND2 i5316 (.O(n7938), .I0(n6_adj_164), .I1(int_Data1[3]));
    AND2 i5494 (.O(n8120), .I0(n8113), .I1(timecnt[11]));
    XOR2 i2_adj_194 (.O(n3758), .I0(n4_adj_17), .I1(n79_adj_111));
    OR2 i6465 (.O(n9108), .I0(int_Data[5]), .I1(n6111));
    AND2 i5501 (.O(n8127), .I0(n8120), .I1(timecnt[12]));
    INV i1150 (.O(n25), .I0(key_out_c_2));
    XOR2 i2_adj_195 (.O(n8399), .I0(n4_adj_177), .I1(n97_adj_49));
    XOR2 i2_adj_196 (.O(n8400), .I0(n4_adj_166), .I1(n73));
    XOR2 i2_adj_197 (.O(n8401), .I0(n4_adj_162), .I1(n49));
    XOR2 i2_adj_198 (.O(n3721), .I0(n4_adj_161), .I1(n124));
    INV i3299 (.O(n4_adj_85), .I0(n5880));
    AND2 i6755 (.O(n9405), .I0(n1298), .I1(n9028));
    INV i3296 (.O(n6_adj_86), .I0(n13));
    OR2 i6756 (.O(n9406), .I0(n9405), .I1(n9404));
    OR2 i6675 (.O(n9325), .I0(n9324), .I1(n9323));
    XOR2 i1_adj_199 (.O(n9035), .I0(n9033), .I1(n7911));
    OR2 i1_adj_200 (.O(n70_adj_57), .I0(n67), .I1(n92));
    AND2 i1_adj_201 (.O(n69), .I0(int_Data1[1]), .I1(n7_adj_89));
    AND2 i6677 (.O(n9327), .I0(n1512), .I1(n9337));
    AND2 i1_adj_202 (.O(n770), .I0(n8964), .I1(n8458));
    OR2 i6678 (.O(led_int_Data0_3__N_59[3]), .I0(n9327), .I1(n9326));
    AND2 i2_adj_203 (.O(n6_adj_99), .I0(n87_adj_109), .I1(n25));
    OR2 i3273 (.O(n5854), .I0(key_in_c_1), .I1(key_in_c_2));
    OR3 i2_adj_204 (.O(n11_adj_115), .I0(n9_adj_47), .I1(key_out_c_3), 
        .I2(n25));
    AND3 i6667 (.O(n9317), .I0(n115), .I1(n29_adj_29), .I2(key_out_c_3));
    OR2 i6623 (.O(n9273), .I0(n9272), .I1(n9271));
    AND2 i3516 (.O(n6111), .I0(n6038), .I1(n6_adj_117));
    OR2 i1786 (.O(n4293), .I0(n1317), .I1(n4292));
    AND2 i6758 (.O(n9408), .I0(n1299), .I1(n539));
    AND2 i1785 (.O(n4292), .I0(n3825), .I1(n5839));
    AND3 i1_adj_205 (.O(n744), .I0(n8464), .I1(n4495), .I2(n8458));
    AND2 i1_adj_206 (.O(n68), .I0(int_Data1[2]), .I1(n7_adj_89));
    INV i6593 (.O(n9243), .I0(n9010));
    OR2 i3616 (.O(n6020), .I0(n6225), .I1(n14_adj_114));
    AND2 i3396 (.O(n3204), .I0(n1511), .I1(n731));
    AND2 i1_adj_207 (.O(n102), .I0(n9316), .I1(n10));
    AND3 i6479 (.O(n9124), .I0(n5953), .I1(n15_adj_106), .I2(n94));
    AND2 i6430 (.O(n9122), .I0(n21_adj_125), .I1(n21));
    INV i3293 (.O(n4_adj_94), .I0(n5874));
    OR2 i6645 (.O(n9295), .I0(n9294), .I1(n9293));
    INV i6588 (.O(n9238), .I0(n15_adj_53));
    INV i6437 (.O(n9_adj_140), .I0(n111));
    INV i3539 (.O(n20), .I0(n6133));
    OR2 i1_adj_208 (.O(n4490), .I0(n4489), .I1(n531));
    OR2 i5570 (.O(n4_adj_183), .I0(n8198), .I1(n8202));
    INV i119 (.O(n101), .I0(n8302));
    OR2 i1_adj_209 (.O(n4491), .I0(n4489), .I1(n563));
    AND2 i1_adj_210 (.O(n8968), .I0(n8467), .I1(n8504));
    XOR2 i1_adj_211 (.O(n8427), .I0(n540), .I1(n8439));
    AND2 i1_adj_212 (.O(led_int_Data1_3__N_385), .I0(n8968), .I1(n8468));
    AND2 i6680 (.O(n9330), .I0(n1512), .I1(n9340));
    OR2 i3499 (.O(n6093), .I0(n6101), .I1(n14));
    OR2 i5617 (.O(n4_adj_76), .I0(n8250), .I1(n8254));
    OR2 i6681 (.O(led_int_Data0_3__N_59[2]), .I0(n9330), .I1(n9329));
    AND2 i5618 (.O(n8254), .I0(n8253), .I1(n3725));
    OR2 i3498 (.O(n862), .I0(n4572), .I1(n796));
    AND2 i5376 (.O(n8001), .I0(n6_adj_171), .I1(n6));
    AND3 i2_adj_213 (.O(n8343), .I0(n6581), .I1(int_Data0[7]), .I2(flag_Data[1]));
    XOR2 i1_adj_214 (.O(n8435), .I0(n12), .I1(int_Data0[6]));
    OR2 i1_adj_215 (.O(n9_adj_47), .I0(key_out_c_1), .I1(key_out_c_0));
    XOR2 i5428 (.O(n78), .I0(n8050), .I1(timecnt[2]));
    OR2 i1738 (.O(n4245), .I0(n1311), .I1(n4244));
    AND2 i1737 (.O(n4244), .I0(n4293), .I1(n5835));
    OR2 i5546 (.O(n8176), .I0(n6_adj_165), .I1(n103));
    AND2 i5508 (.O(n8134), .I0(n8127), .I1(timecnt[13]));
    XOR2 i1_adj_216 (.O(n8506), .I0(n5955), .I1(n8425));
    AND2 i3238 (.O(n93), .I0(n29), .I1(n76_adj_12));
    OR2 i3528 (.O(n6123), .I0(n8_adj_15), .I1(int_Data[1]));
    INV i6433 (.O(n8986), .I0(n9072));
    INV i6636 (.O(n9286), .I0(n9118));
    AND2 i5438 (.O(n8064), .I0(n8057), .I1(timecnt[3]));
    AND2 i6683 (.O(n9333), .I0(n1512), .I1(n9343));
    AND2 i6616 (.O(n9266), .I0(n1464), .I1(n3830));
    AND3 i6664 (.O(n9314), .I0(n4_adj_85), .I1(n31), .I2(n99));
    AND2 i6760 (.O(n9410), .I0(n8354), .I1(n9409));
    AND2 i6757 (.O(n9407), .I0(n4491), .I1(n9364));
    AND2 i6754 (.O(n9404), .I0(n8354), .I1(n9403));
    AND2 i6751 (.O(n9401), .I0(n4491), .I1(n9361));
    AND3 i6661 (.O(n9311), .I0(n4540), .I1(n29_adj_29), .I2(n25));
    AND2 i6748 (.O(n9398), .I0(n8354), .I1(n9397));
    AND2 i6745 (.O(n9395), .I0(n4491), .I1(n9358));
    AND2 i6742 (.O(n9392), .I0(n8354), .I1(n9391));
    AND2 i6739 (.O(n9389), .I0(n4491), .I1(n9355));
    AND2 i6736 (.O(n9386), .I0(n8354), .I1(n9385));
    AND2 i6733 (.O(n9383), .I0(n4491), .I1(n9352));
    INV i1927 (.O(n1488), .I0(n4462));
    XOR2 i2_adj_217 (.O(n9_adj_56), .I0(n10_adj_174), .I1(n169));
    XOR2 i1_adj_218 (.O(n4_adj_139), .I0(int_Data[3]), .I1(n3204));
    AND4 i6658 (.O(n9308), .I0(key_in_c_3), .I1(key_out_c_3), .I2(n31), 
         .I3(n6_adj_24));
    AND2 i6730 (.O(n9380), .I0(n8354), .I1(n9379));
    OR2 i1_adj_219 (.O(n24), .I0(n41_adj_154), .I1(n28_adj_122));
    AND2 i6727 (.O(n9377), .I0(n4491), .I1(n9349));
    AND2 i6724 (.O(n9374), .I0(n8354), .I1(n9373));
    XOR2 i1_adj_220 (.O(n4471), .I0(n6368), .I1(n8433));
    AND2 i5571 (.O(n8202), .I0(n8201), .I1(n3760));
    AND2 i6472 (.O(n9116), .I0(n8988), .I1(n6123));
    OR2 i5547 (.O(n8_adj_167), .I0(n8173), .I1(n8177));
    OR2 i6432 (.O(n9072), .I0(flag_Cal[0]), .I1(flag_Cal[1]));
    OR2 i5369 (.O(n7995), .I0(n4_adj_129), .I1(n7_adj_13));
    OR2 i1_adj_221 (.O(n49_adj_150), .I0(n28_adj_151), .I1(n4554));
    OR2 i5370 (.O(n6_adj_171), .I0(n7992), .I1(n7996));
    XOR2 i1_adj_222 (.O(n8441), .I0(n8_adj_172), .I1(int_Data0[4]));
    AND2 i1_adj_223 (.O(n67), .I0(int_Data1[0]), .I1(n7_adj_89));
    AND2 i3497 (.O(led_int_Data1_3__N_63[2]), .I0(n6089), .I1(n862));
    OR2 i1_adj_224 (.O(n4_adj_64), .I0(n31), .I1(key_in_c_1));
    AND2 i1_adj_225 (.O(n9002), .I0(n8982), .I1(n6093));
    INV i1244 (.O(n20_adj_1), .I0(key_out_c_0));
    OR2 i3277 (.O(n1556), .I0(n5797), .I1(int_Data[2]));
    XOR2 i3_adj_226 (.O(n10_adj_3), .I0(n8_adj_167), .I1(n148));
    XOR2 i4_adj_227 (.O(n11), .I0(n8_adj_77), .I1(n127));
    AND2 i1_adj_228 (.O(n8345), .I0(n5797), .I1(int_Data[2]));
    AND3 i6655 (.O(n9305), .I0(n84), .I1(n10), .I2(key_in_c_0));
    AND2 i6652 (.O(n9302), .I0(n5869), .I1(n9412));
    OR2 i1_adj_229 (.O(n9022), .I0(n22_adj_19), .I1(flag_Data[0]));
    AND2 i3241 (.O(n94_adj_72), .I0(n29), .I1(n77));
    AND2 i1656 (.O(n4149), .I0(n4148), .I1(int_Data[2]));
    AND2 i3380 (.O(led_int_Data1_3__N_63[1]), .I0(n1511), .I1(led_int_Data1_3__N_381[1]));
    OR2 i6684 (.O(led_int_Data0_3__N_59[1]), .I0(n9333), .I1(n9332));
    OR2 i3490 (.O(led_int_Data1_3__N_381[1]), .I0(n4_adj_157), .I1(n8744));
    AND2 i1_adj_230 (.O(n8993), .I0(n8991), .I1(n5913));
    OR2 i3737 (.O(n6368), .I0(n6314), .I1(n534));
    OR2 i5377 (.O(n8004), .I0(n6_adj_171), .I1(n6));
    AND2 i6649 (.O(n9299), .I0(n5869), .I1(n9406));
    OR2 i1_adj_231 (.O(n4495), .I0(n4492), .I1(n4535));
    AND2 i1627 (.O(n4_adj_14), .I0(int_Data[1]), .I1(n4355));
    AND2 i6686 (.O(n9336), .I0(n757), .I1(n7_adj_136));
    AND3 i1_adj_232 (.O(n8971), .I0(key_out_c_3), .I1(n15_adj_81), .I2(key_in_c_0));
    AND2 i1_adj_233 (.O(n4_adj_184), .I0(n8498), .I1(n10_adj_18));
    AND2 i1_adj_234 (.O(n4535), .I0(n6038), .I1(n6_adj_137));
    AND3 i6556 (.O(n9205), .I0(n8982), .I1(n5913), .I2(n6150));
    OR2 i1604 (.O(n3825), .I0(n1323), .I1(n4090));
    AND4 i6646 (.O(n9296), .I0(key_out_c_0), .I1(n10), .I2(n25), .I3(key_in_c_2));
    AND2 i1603 (.O(n4090), .I0(n1329), .I1(n5843));
    AND2 i1_adj_235 (.O(n41_adj_154), .I0(n40), .I1(n21_adj_132));
    AND2 i5548 (.O(n8177), .I0(n8176), .I1(n82_adj_60));
    XOR2 i1_adj_236 (.O(n4473), .I0(n6314), .I1(n8435));
    XOR2 i104 (.O(n92_adj_147), .I0(key_out_c_3), .I1(key_out_c_0));
    OR2 i3538 (.O(n6133), .I0(n5874), .I1(key_out_c_0));
    AND2 i6643 (.O(n9293), .I0(n5869), .I1(n9400));
    XOR2 i1_adj_237 (.O(n4_adj_191), .I0(n6_adj_182), .I1(n3758));
    OR2 i1585 (.O(n4067), .I0(n1305), .I1(n4066));
    OR2 i1_adj_238 (.O(n68_adj_145), .I0(n8310), .I1(n4_adj_68));
    AND2 i1_adj_239 (.O(n28_adj_122), .I0(n15_adj_73), .I1(n14_adj_83));
    AND2 i1584 (.O(n4066), .I0(n4245), .I1(n9006));
    INV i1146 (.O(n19), .I0(key_out_c_1));
    AND2 i5424 (.O(n8050), .I0(timecnt[0]), .I1(timecnt[1]));
    XOR2 i5 (.O(n12_adj_199), .I0(n10_adj_3), .I1(n9_adj_56));
    XOR2 i2_adj_240 (.O(n4459), .I0(n4_adj_158), .I1(n4_adj_14));
    OR2 i6687 (.O(n9337), .I0(n9336), .I1(n9335));
    AND2 i1_adj_241 (.O(n4540), .I0(key_out_c_1), .I1(key_in_c_2));
    XOR2 i48 (.O(n50), .I0(key_in_c_1), .I1(key_in_c_0));
    AND2 i6689 (.O(n9339), .I0(n757), .I1(int_Data[2]));
    OR2 i1_adj_242 (.O(n4_adj_157), .I0(n744), .I1(n731));
    AND2 i1_adj_243 (.O(n4587), .I0(n4586), .I1(int_Data0_7__N_151[2]));
    XOR2 i49 (.O(n34_adj_144), .I0(key_out_c_2), .I1(key_out_c_1));
    AND3 i2_adj_244 (.O(n8348), .I0(n4789), .I1(int_Data0[4]), .I2(flag_Data[1]));
    INV i5419 (.O(n80), .I0(timecnt[0]));
    AND2 i1_adj_245 (.O(n82_adj_51), .I0(n3842), .I1(flag_Data[0]));
    OR2 i1_adj_246 (.O(n4561), .I0(int_Data[6]), .I1(int_Data[7]));
    OR2 i1_adj_247 (.O(n4492), .I0(n4561), .I1(int_Data[5]));
    OR2 i1_adj_248 (.O(n4564), .I0(n4561), .I1(n8326));
    OR2 i3544 (.O(n5883), .I0(n6141), .I1(n11_adj_7));
    OR2 i1_adj_249 (.O(n4_adj_195), .I0(key_in_c_0), .I1(n10));
    OR3 i1_adj_250 (.O(n4567), .I0(n10_adj_79), .I1(int_Data[5]), .I2(n6_adj_137));
    OR2 i1535 (.O(n6_adj_187), .I0(key_out_c_2), .I1(n7_adj_89));
    INV equal_22_i8 (.O(n92), .I0(n14_adj_20));
    INV i2163 (.O(n9_adj_27), .I0(key_in_c_2));
    INV i3305 (.O(n5887), .I0(n3967));
    XOR2 i2_adj_251 (.O(n8398), .I0(n4_adj_149), .I1(n121));
    INV i3274 (.O(n5_adj_93), .I0(n5854));
    OR2 i1_adj_252 (.O(n40), .I0(n12_adj_138), .I1(n18));
    INV i6533 (.O(n9051), .I0(n9180));
    OR2 i3298 (.O(n5880), .I0(key_out_c_0), .I1(key_out_c_3));
    INV i78 (.O(n78_adj_33), .I0(flag_Cal[0]));
    INV i3740 (.O(n4787), .I0(n9003));
    XOR2 i2_adj_253 (.O(n3759), .I0(n4_adj_141), .I1(n55_adj_134));
    INV i6562 (.O(n9016), .I0(n9211));
    XOR2 i52 (.O(n38_adj_142), .I0(key_in_c_3), .I1(key_in_c_2));
    OR2 equal_412_i14 (.O(n14_adj_20), .I0(n3842), .I1(flag_Data[0]));
    INV i3215 (.O(n1207), .I0(n5795));
    AND2 i6474 (.O(n9118), .I0(n8354), .I1(n4489));
    AND2 i5623 (.O(n8259), .I0(n4_adj_76), .I1(n73));
    OR2 i3292 (.O(n5874), .I0(key_out_c_2), .I1(key_out_c_1));
    AND3 i2_adj_254 (.O(n8300), .I0(n101), .I1(int_Data1[3]), .I2(n5887));
    AND2 i1_adj_255 (.O(n66), .I0(int_Data1[3]), .I1(n7_adj_89));
    OR2 i2_adj_256 (.O(n24_adj_189), .I0(n4_adj_135), .I1(n13));
    OR2 i6690 (.O(n9340), .I0(n9339), .I1(n9338));
    OR2 i1_adj_257 (.O(n4639), .I0(n4638), .I1(n8340));
    AND4 i6625 (.O(n9275), .I0(n6_adj_98), .I1(n97_adj_28), .I2(key_in_c_0), 
         .I3(n9_adj_27));
    OR2 i1_adj_258 (.O(n4645), .I0(n4644), .I1(n8339));
    OR3 i2_adj_259 (.O(n4681), .I0(n1208), .I1(n7_adj_89), .I2(n1207));
    AND2 mult_119_i2 (.O(n7911), .I0(int_Data1[0]), .I1(int_Data0[0]));
    AND2 mult_119_i4 (.O(n5), .I0(int_Data1[1]), .I1(int_Data0[0]));
    AND2 mult_119_i6 (.O(n8_adj_38), .I0(int_Data1[2]), .I1(int_Data0[0]));
    AND2 mult_119_i8 (.O(n11_adj_155), .I0(int_Data1[3]), .I1(int_Data0[0]));
    AND2 i3679 (.O(n9_adj_160), .I0(n5999), .I1(n5843));
    AND2 mult_119_i18 (.O(n25_adj_159), .I0(int_Data1[0]), .I1(int_Data0[1]));
    AND2 mult_119_i20 (.O(n28_adj_5), .I0(int_Data1[1]), .I1(int_Data0[1]));
    AND2 i6692 (.O(n9342), .I0(n757), .I1(int_Data[1]));
    AND2 mult_119_i22 (.O(n31_adj_50), .I0(int_Data1[2]), .I1(int_Data0[1]));
    OR2 i6693 (.O(n9343), .I0(n9342), .I1(n9341));
    AND2 mult_119_i24 (.O(n34), .I0(int_Data1[3]), .I1(int_Data0[1]));
    OR2 i3551 (.O(n6150), .I0(n6225), .I1(n14_adj_107));
    AND2 mult_119_i34 (.O(n49), .I0(int_Data1[0]), .I1(int_Data0[2]));
    INV i3267 (.O(n4_adj_100), .I0(n10_adj_121));
    INV i3265 (.O(n1329), .I0(n5999));
    INV i5798 (.O(n535), .I0(n8437));
    INV i3261 (.O(n1323), .I0(n5841));
    AND2 mult_119_i36 (.O(n52), .I0(int_Data1[1]), .I1(int_Data0[2]));
    AND2 mult_119_i38 (.O(n55_adj_134), .I0(int_Data1[2]), .I1(int_Data0[2]));
    OR2 i1_adj_260 (.O(n3967), .I0(n92), .I1(n82_adj_51));
    AND2 i6640 (.O(n9290), .I0(n3842), .I1(led_int_Data2_3__N_111[1]));
    AND2 mult_119_i40 (.O(n58), .I0(int_Data1[3]), .I1(int_Data0[2]));
    OR2 i5317 (.O(n7941), .I0(n6_adj_164), .I1(int_Data1[3]));
    AND2 mult_119_i50 (.O(n73), .I0(int_Data1[0]), .I1(int_Data0[3]));
    AND2 mult_119_i52 (.O(n76), .I0(int_Data1[1]), .I1(int_Data0[3]));
    AND2 mult_119_i54 (.O(n79_adj_111), .I0(int_Data1[2]), .I1(int_Data0[3]));
    AND2 mult_119_i56 (.O(n82_adj_60), .I0(int_Data1[3]), .I1(int_Data0[3]));
    AND2 mult_119_i66 (.O(n97_adj_49), .I0(int_Data1[0]), .I1(int_Data0[4]));
    AND2 mult_119_i68 (.O(n100_adj_128), .I0(int_Data1[1]), .I1(int_Data0[4]));
    OR2 i5318 (.O(n8_adj_173), .I0(n7938), .I1(n7942));
    AND2 mult_119_i70 (.O(n103), .I0(int_Data1[2]), .I1(int_Data0[4]));
    GND i1 (.X(n929));
    INV i3257 (.O(n1317), .I0(n5837));
    AND2 i6587 (.O(n13_adj_41), .I0(n9273), .I1(n9236));
    AND2 mult_119_i72 (.O(n106), .I0(int_Data1[3]), .I1(int_Data0[4]));
    OR2 i6478 (.O(n9123), .I0(n9122), .I1(n19_adj_148));
    AND2 mult_119_i82 (.O(n121), .I0(int_Data1[0]), .I1(int_Data0[5]));
    AND2 mult_119_i84 (.O(n124), .I0(int_Data1[1]), .I1(int_Data0[5]));
    AND3 i2_adj_261 (.O(n8315), .I0(n9_adj_27), .I1(key_in_c_1), .I2(n6_adj_99));
    INV i3253 (.O(n1311), .I0(n9007));
    
endmodule
//
// Verilog Description of module AND2
// module not written out since it is a black-box. 
//

//
// Verilog Description of module AND5
// module not written out since it is a black-box. 
//

//
// Verilog Description of module OR2
// module not written out since it is a black-box. 
//

//
// Verilog Description of module XOR2
// module not written out since it is a black-box. 
//

//
// Verilog Description of module INV
// module not written out since it is a black-box. 
//

//
// Verilog Description of module AND3
// module not written out since it is a black-box. 
//

//
// Verilog Description of module AND4
// module not written out since it is a black-box. 
//

//
// Verilog Description of module OR3
// module not written out since it is a black-box. 
//

//
// Verilog Description of module OR5
// module not written out since it is a black-box. 
//

//
// Verilog Description of module AND6
// module not written out since it is a black-box. 
//

//
// Verilog Description of module OR4
// module not written out since it is a black-box. 
//

//
// Verilog Description of module VCC
// module not written out since it is a black-box. 
//

//
// Verilog Description of module OR6
// module not written out since it is a black-box. 
//

//
// Verilog Description of module GND
// module not written out since it is a black-box. 
//

