module musicplayer(reset,clk,Clock4Hz,EnSp);
input reset; 
input  clk;
input  Clock4Hz;
output EnSp;

reg tone,origin,CntSp,sp,EnSp;
reg [7:0] led;
reg [7:0] CntSone;
always@(tone,reset)
begin
     if(reset==0)
    begin
    EnSp<=0; //EnSp?????????????????0?????
    led<=8'b11111111;//LED ?????
    end
    else
        begin
            case(tone)//tone????????????
               0:begin led<=8'b11111111;EnSp<=0;end//???????
               1:begin origin<=11468; led<=8'b11111110; EnSp<=1;end //???? 1
               2:begin origin<=10215; led<=8'b11111100; EnSp<=1; end //???? 2
               3:begin origin<=9099;led<=8'b11111000;EnSp<=1;end//????3
               4:begin origin<=8591; led<=8'b11110000; EnSp<=1; end //???? 4
               5:begin origin<=7653; led<=8'b11100000; EnSp<=1; end //???? 5
               6:begin origin<=6818; led<=8'b11000000; EnSp<=1; end //???? 6
               7:begin origin<=6074;led<=8'b10000000;EnSp<=1;end//????7
               8:begin origin<=5733; led<=8'b00000000; EnSp<=1; end //????
               default:begin led<=8'b11111111; EnSp<=0;end //???????
            endcase
        end
end

always@(posedge clk or negedge reset) //clk ?????6MHz
begin
    if(reset==0)
        begin
           CntSp<=0;//CntSp????????????????????????
           sp<=1; //sp ?????????????????????
        end
    else if(EnSp==1)
    //origin???????????????sp?????????????????????????????
    //origin ???????????????sp ????????????????????????????
	    begin
           if(CntSp==0) begin CntSp<=origin; sp<=~sp; end
           else CntSp<=CntSp-1;
        end
    else sp<=1;
end

//????
//?????????????????????????�??????????????????
//???????????????????
always@(posedge Clock4Hz or negedge reset) //Clock4Hz?4Hz??????????????????????
begin
     if(reset==0) CntSone<=0;//CntSone????????????????
     else
          begin
             case(CntSone)
                  0: tone<=1;
                  2: tone<=1;
                  4: tone<=5;
                  6: tone<=5;
				  8: tone<=6;
				  10: tone<=6;
                  12: tone<=5;
                  13: tone<=5;
				  
                  16: tone<=4;
				  18: tone<=4;
                  20: tone<=3;
                  22: tone<=3;
                  24: tone<=2;
				  26: tone<=2;
                  28: tone<=1;
                  29: tone<=1;
				  
				  32: tone<=5;
				  34: tone<=5;
                  36: tone<=4;
                  38: tone<=4;
                  40: tone<=3;
				  42: tone<=3;
                  44: tone<=2;
                  45: tone<=2;
				  
				  48: tone<=5;
				  50: tone<=5;
                  52: tone<=4;
                  54: tone<=4;
                  56: tone<=3;
				  58: tone<=3;
                  60: tone<=2;
                  61: tone<=2;
                  
                  default: tone<=0;
             endcase
             if(CntSone==67) CntSone<=0;
             else CntSone<=CntSone+1;
          end
end
endmodule