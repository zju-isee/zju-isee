module DISPLAY(clk,reset,num1,num2,num3,num4,LED_A,LED_B,LED_C,LED_D,LED_E,LED_F,LED_G,LED_VCC1,LED_VCC2,LED_VCC3,LED_VCC4);
input clk;                      //ʱ���ź�
input reset;                    //��λ�ź�
input [3:0] num1;             //���������
input [3:0] num2;             //���������
input [3:0] num3;             //���������
input [3:0] num4;             //���������

output reg LED_A,LED_B,LED_C,LED_D,LED_E,LED_F,LED_G,LED_VCC1,LED_VCC2,LED_VCC3,LED_VCC4;

reg [1:0] scancnt;
reg [12:0] count;



always @(posedge clk or negedge reset)
begin
    if(reset==1'b0)count=0;
    else if(count==5999)
        begin
            count=0;
            if(scancnt==3)scancnt=0;
            else scancnt=scancnt+1;
        end
    else count=count+1;
end

always @(posedge clk) begin
    if(reset==1'b0)
        begin
            LED_A=1;LED_B=1;LED_C=1;LED_D=1;
            LED_E=1;LED_F=1;LED_G=1;//�߶���
            LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
            LED_VCC4=0;//ǧ��ʮ��λ
        end
    else if(scancnt==0)
        begin
            case (num1)
                0:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=0;
                    LED_E=0;LED_F=0;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=1;//ǧ��ʮ��λ
                end
                1:begin
                    LED_A=1;LED_B=0;LED_C=0;LED_D=1;
                    LED_E=1;LED_F=1;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=1;//ǧ��ʮ��λ
                end
                2:begin
                    LED_A=0;LED_B=0;LED_C=1;LED_D=0;
                    LED_E=0;LED_F=1;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=1;//ǧ��ʮ��λ
                end
                3:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=0;
                    LED_E=1;LED_F=1;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=1;//ǧ��ʮ��λ
                end
                4:begin
                    LED_A=1;LED_B=0;LED_C=0;LED_D=1;
                    LED_E=1;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=1;//ǧ��ʮ��λ
                end
                5:begin
                    LED_A=0;LED_B=1;LED_C=0;LED_D=0;
                    LED_E=1;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=1;//ǧ��ʮ��λ
                end
                6:begin
                    LED_A=0;LED_B=1;LED_C=0;LED_D=0;
                    LED_E=0;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=1;//ǧ��ʮ��λ
                    end
                7:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=1;
                    LED_E=1;LED_F=1;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=1;//ǧ��ʮ��λ
                end
                8:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=0;
                    LED_E=0;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=1;//ǧ��ʮ��λ 
                end
                9:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=0;
                    LED_E=1;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=1;//ǧ��ʮ��λ
                end
                10:begin
                    LED_A=1;LED_B=1;LED_C=1;LED_D=1;
                    LED_E=1;LED_F=1;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=1;//ǧ��ʮ��λ
                end 
                default:begin
                    LED_A=1;LED_B=1;LED_C=1;LED_D=1;
                    LED_E=1;LED_F=1;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=1;//ǧ��ʮ��λ
                end
            endcase
        end
    else if(scancnt==1)
        begin
            case (num2)
                0:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=0;
                    LED_E=0;LED_F=0;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=1;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                1:begin
                    LED_A=1;LED_B=0;LED_C=0;LED_D=1;
                    LED_E=1;LED_F=1;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=1;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                2:begin
                    LED_A=0;LED_B=0;LED_C=1;LED_D=0;
                    LED_E=0;LED_F=1;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=1;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                3:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=0;
                    LED_E=1;LED_F=1;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=1;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                4:begin
                    LED_A=1;LED_B=0;LED_C=0;LED_D=1;
                    LED_E=1;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=1;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                5:begin
                    LED_A=0;LED_B=1;LED_C=0;LED_D=0;
                    LED_E=1;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=1;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                6:begin
                    LED_A=0;LED_B=1;LED_C=0;LED_D=0;
                    LED_E=0;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=1;
                    LED_VCC4=0;//ǧ��ʮ��λ
                    end
                7:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=1;
                    LED_E=1;LED_F=1;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=1;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                8:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=0;
                    LED_E=0;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=1;
                    LED_VCC4=0;//ǧ��ʮ��λ 
                end
                9:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=0;
                    LED_E=1;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=1;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                10:begin
                    LED_A=1;LED_B=1;LED_C=1;LED_D=1;
                    LED_E=1;LED_F=1;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=1;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                default:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=0;
                    LED_E=0;LED_F=0;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=1;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
            endcase
        end
    else if(scancnt==2)
        begin
            case (num3)
                0:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=0;
                    LED_E=0;LED_F=0;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=1;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                1:begin
                    LED_A=1;LED_B=0;LED_C=0;LED_D=1;
                    LED_E=1;LED_F=1;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=1;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                2:begin
                    LED_A=0;LED_B=0;LED_C=1;LED_D=0;
                    LED_E=0;LED_F=1;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=1;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                3:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=0;
                    LED_E=1;LED_F=1;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=1;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                4:begin
                    LED_A=1;LED_B=0;LED_C=0;LED_D=1;
                    LED_E=1;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=1;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                5:begin
                    LED_A=0;LED_B=1;LED_C=0;LED_D=0;
                    LED_E=1;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=1;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                6:begin
                    LED_A=0;LED_B=1;LED_C=0;LED_D=0;
                    LED_E=0;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=1;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                    end
                7:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=1;
                    LED_E=1;LED_F=1;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=1;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                8:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=0;
                    LED_E=0;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=1;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ 
                end
                9:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=0;
                    LED_E=1;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=1;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                10:begin
                    LED_A=1;LED_B=1;LED_C=1;LED_D=1;
                    LED_E=1;LED_F=1;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=1;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                11:begin
                    LED_A=1;LED_B=1;LED_C=1;LED_D=1;
                    LED_E=1;LED_F=1;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=1;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                default:begin
                    LED_A=1;LED_B=1;LED_C=1;LED_D=1;
                    LED_E=1;LED_F=1;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=1;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
            endcase
        end
    else if(scancnt==3)
        begin
            case (num4)
                0:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=0;
                    LED_E=0;LED_F=0;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                1:begin
                    LED_A=1;LED_B=0;LED_C=0;LED_D=1;
                    LED_E=1;LED_F=1;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                2:begin
                    LED_A=0;LED_B=0;LED_C=1;LED_D=0;
                    LED_E=0;LED_F=1;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                3:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=0;
                    LED_E=1;LED_F=1;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                4:begin
                    LED_A=1;LED_B=0;LED_C=0;LED_D=1;
                    LED_E=1;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                5:begin
                    LED_A=0;LED_B=1;LED_C=0;LED_D=0;
                    LED_E=1;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                6:begin
                    LED_A=0;LED_B=1;LED_C=0;LED_D=0;
                    LED_E=0;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                    end
                7:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=1;
                    LED_E=1;LED_F=1;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                8:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=0;
                    LED_E=0;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ 
                end
                9:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=0;
                    LED_E=1;LED_F=0;LED_G=0;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
                default:begin
                    LED_A=0;LED_B=0;LED_C=0;LED_D=0;
                    LED_E=0;LED_F=0;LED_G=1;//�߶���
                    LED_VCC1=0;LED_VCC2=0;LED_VCC3=0;
                    LED_VCC4=0;//ǧ��ʮ��λ
                end
            endcase
        end
    end
endmodule

